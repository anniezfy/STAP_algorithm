module CORDIC_CR_ORIGIN(
  input         clock,
  input         reset,
  input  [63:0] io_x,
  input  [63:0] io_y,
  input  [63:0] io_theta,
  output [63:0] io_x_n,
  output [63:0] io_y_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] current_x_0; // @[Cordic_CR.scala 42:43]
  reg [63:0] current_x_1; // @[Cordic_CR.scala 42:43]
  reg [63:0] current_x_2; // @[Cordic_CR.scala 42:43]
  reg [63:0] current_x_3; // @[Cordic_CR.scala 42:43]
  reg [63:0] current_x_4; // @[Cordic_CR.scala 42:43]
  reg [63:0] current_x_5; // @[Cordic_CR.scala 42:43]
  reg [63:0] current_x_6; // @[Cordic_CR.scala 42:43]
  reg [63:0] current_x_7; // @[Cordic_CR.scala 42:43]
  reg [63:0] current_x_8; // @[Cordic_CR.scala 42:43]
  reg [63:0] current_x_9; // @[Cordic_CR.scala 42:43]
  reg [63:0] current_x_10; // @[Cordic_CR.scala 42:43]
  reg [63:0] current_x_11; // @[Cordic_CR.scala 42:43]
  reg [63:0] current_x_12; // @[Cordic_CR.scala 42:43]
  reg [63:0] current_x_13; // @[Cordic_CR.scala 42:43]
  reg [63:0] current_x_14; // @[Cordic_CR.scala 42:43]
  reg [63:0] current_y_0; // @[Cordic_CR.scala 43:43]
  reg [63:0] current_y_1; // @[Cordic_CR.scala 43:43]
  reg [63:0] current_y_2; // @[Cordic_CR.scala 43:43]
  reg [63:0] current_y_3; // @[Cordic_CR.scala 43:43]
  reg [63:0] current_y_4; // @[Cordic_CR.scala 43:43]
  reg [63:0] current_y_5; // @[Cordic_CR.scala 43:43]
  reg [63:0] current_y_6; // @[Cordic_CR.scala 43:43]
  reg [63:0] current_y_7; // @[Cordic_CR.scala 43:43]
  reg [63:0] current_y_8; // @[Cordic_CR.scala 43:43]
  reg [63:0] current_y_9; // @[Cordic_CR.scala 43:43]
  reg [63:0] current_y_10; // @[Cordic_CR.scala 43:43]
  reg [63:0] current_y_11; // @[Cordic_CR.scala 43:43]
  reg [63:0] current_y_12; // @[Cordic_CR.scala 43:43]
  reg [63:0] current_y_13; // @[Cordic_CR.scala 43:43]
  reg [63:0] current_y_14; // @[Cordic_CR.scala 43:43]
  reg [63:0] current_theta_0; // @[Cordic_CR.scala 44:47]
  reg [63:0] current_theta_1; // @[Cordic_CR.scala 44:47]
  reg [63:0] current_theta_2; // @[Cordic_CR.scala 44:47]
  reg [63:0] current_theta_3; // @[Cordic_CR.scala 44:47]
  reg [63:0] current_theta_4; // @[Cordic_CR.scala 44:47]
  reg [63:0] current_theta_5; // @[Cordic_CR.scala 44:47]
  reg [63:0] current_theta_6; // @[Cordic_CR.scala 44:47]
  reg [63:0] current_theta_7; // @[Cordic_CR.scala 44:47]
  reg [63:0] current_theta_8; // @[Cordic_CR.scala 44:47]
  reg [63:0] current_theta_9; // @[Cordic_CR.scala 44:47]
  reg [63:0] current_theta_10; // @[Cordic_CR.scala 44:47]
  reg [63:0] current_theta_11; // @[Cordic_CR.scala 44:47]
  reg [63:0] current_theta_12; // @[Cordic_CR.scala 44:47]
  reg [63:0] current_theta_13; // @[Cordic_CR.scala 44:47]
  wire [63:0] _current_x_0_T_2 = $signed(io_x) + $signed(io_y); // @[Cordic_CR.scala 54:30]
  wire [63:0] _current_y_0_T_2 = 64'sh0 - $signed(io_x); // @[Cordic_CR.scala 55:25]
  wire [63:0] _current_y_0_T_5 = $signed(_current_y_0_T_2) + $signed(io_y); // @[Cordic_CR.scala 55:31]
  wire [63:0] _current_theta_0_T_2 = $signed(io_theta) + 64'sh2d00000000; // @[Cordic_CR.scala 56:38]
  wire [63:0] _current_x_0_T_5 = $signed(io_x) - $signed(io_y); // @[Cordic_CR.scala 58:30]
  wire [63:0] _current_theta_0_T_5 = $signed(io_theta) - 64'sh2d00000000; // @[Cordic_CR.scala 60:38]
  wire [62:0] _current_x_1_T = current_y_0[63:1]; // @[Cordic_CR.scala 64:62]
  wire [63:0] _GEN_45 = {{1{_current_x_1_T[62]}},_current_x_1_T}; // @[Cordic_CR.scala 64:42]
  wire [63:0] _current_x_1_T_3 = $signed(current_x_0) + $signed(_GEN_45); // @[Cordic_CR.scala 64:42]
  wire [62:0] _current_y_1_T = current_x_0[63:1]; // @[Cordic_CR.scala 65:62]
  wire [63:0] _GEN_46 = {{1{_current_y_1_T[62]}},_current_y_1_T}; // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_y_1_T_3 = $signed(current_y_0) - $signed(_GEN_46); // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_theta_1_T_2 = $signed(current_theta_0) + 64'sh1a90a731a6; // @[Cordic_CR.scala 66:50]
  wire [63:0] _current_x_1_T_7 = $signed(current_x_0) - $signed(_GEN_45); // @[Cordic_CR.scala 68:42]
  wire [63:0] _current_y_1_T_7 = $signed(current_y_0) + $signed(_GEN_46); // @[Cordic_CR.scala 69:42]
  wire [63:0] _current_theta_1_T_5 = $signed(current_theta_0) - 64'sh1a90a731a6; // @[Cordic_CR.scala 70:50]
  wire [61:0] _current_x_2_T = current_y_1[63:2]; // @[Cordic_CR.scala 64:62]
  wire [63:0] _GEN_49 = {{2{_current_x_2_T[61]}},_current_x_2_T}; // @[Cordic_CR.scala 64:42]
  wire [63:0] _current_x_2_T_3 = $signed(current_x_1) + $signed(_GEN_49); // @[Cordic_CR.scala 64:42]
  wire [61:0] _current_y_2_T = current_x_1[63:2]; // @[Cordic_CR.scala 65:62]
  wire [63:0] _GEN_50 = {{2{_current_y_2_T[61]}},_current_y_2_T}; // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_y_2_T_3 = $signed(current_y_1) - $signed(_GEN_50); // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_theta_2_T_2 = $signed(current_theta_1) + 64'she0947407d; // @[Cordic_CR.scala 66:50]
  wire [63:0] _current_x_2_T_7 = $signed(current_x_1) - $signed(_GEN_49); // @[Cordic_CR.scala 68:42]
  wire [63:0] _current_y_2_T_7 = $signed(current_y_1) + $signed(_GEN_50); // @[Cordic_CR.scala 69:42]
  wire [63:0] _current_theta_2_T_5 = $signed(current_theta_1) - 64'she0947407d; // @[Cordic_CR.scala 70:50]
  wire [60:0] _current_x_3_T = current_y_2[63:3]; // @[Cordic_CR.scala 64:62]
  wire [63:0] _GEN_53 = {{3{_current_x_3_T[60]}},_current_x_3_T}; // @[Cordic_CR.scala 64:42]
  wire [63:0] _current_x_3_T_3 = $signed(current_x_2) + $signed(_GEN_53); // @[Cordic_CR.scala 64:42]
  wire [60:0] _current_y_3_T = current_x_2[63:3]; // @[Cordic_CR.scala 65:62]
  wire [63:0] _GEN_54 = {{3{_current_y_3_T[60]}},_current_y_3_T}; // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_y_3_T_3 = $signed(current_y_2) - $signed(_GEN_54); // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_theta_3_T_2 = $signed(current_theta_2) + 64'sh72001124a; // @[Cordic_CR.scala 66:50]
  wire [63:0] _current_x_3_T_7 = $signed(current_x_2) - $signed(_GEN_53); // @[Cordic_CR.scala 68:42]
  wire [63:0] _current_y_3_T_7 = $signed(current_y_2) + $signed(_GEN_54); // @[Cordic_CR.scala 69:42]
  wire [63:0] _current_theta_3_T_5 = $signed(current_theta_2) - 64'sh72001124a; // @[Cordic_CR.scala 70:50]
  wire [59:0] _current_x_4_T = current_y_3[63:4]; // @[Cordic_CR.scala 64:62]
  wire [63:0] _GEN_57 = {{4{_current_x_4_T[59]}},_current_x_4_T}; // @[Cordic_CR.scala 64:42]
  wire [63:0] _current_x_4_T_3 = $signed(current_x_3) + $signed(_GEN_57); // @[Cordic_CR.scala 64:42]
  wire [59:0] _current_y_4_T = current_x_3[63:4]; // @[Cordic_CR.scala 65:62]
  wire [63:0] _GEN_58 = {{4{_current_y_4_T[59]}},_current_y_4_T}; // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_y_4_T_3 = $signed(current_y_3) - $signed(_GEN_58); // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_theta_4_T_2 = $signed(current_theta_3) + 64'sh3938aa64c; // @[Cordic_CR.scala 66:50]
  wire [63:0] _current_x_4_T_7 = $signed(current_x_3) - $signed(_GEN_57); // @[Cordic_CR.scala 68:42]
  wire [63:0] _current_y_4_T_7 = $signed(current_y_3) + $signed(_GEN_58); // @[Cordic_CR.scala 69:42]
  wire [63:0] _current_theta_4_T_5 = $signed(current_theta_3) - 64'sh3938aa64c; // @[Cordic_CR.scala 70:50]
  wire [58:0] _current_x_5_T = current_y_4[63:5]; // @[Cordic_CR.scala 64:62]
  wire [63:0] _GEN_61 = {{5{_current_x_5_T[58]}},_current_x_5_T}; // @[Cordic_CR.scala 64:42]
  wire [63:0] _current_x_5_T_3 = $signed(current_x_4) + $signed(_GEN_61); // @[Cordic_CR.scala 64:42]
  wire [58:0] _current_y_5_T = current_x_4[63:5]; // @[Cordic_CR.scala 65:62]
  wire [63:0] _GEN_62 = {{5{_current_y_5_T[58]}},_current_y_5_T}; // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_y_5_T_3 = $signed(current_y_4) - $signed(_GEN_62); // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_theta_5_T_2 = $signed(current_theta_4) + 64'sh1ca3794e5; // @[Cordic_CR.scala 66:50]
  wire [63:0] _current_x_5_T_7 = $signed(current_x_4) - $signed(_GEN_61); // @[Cordic_CR.scala 68:42]
  wire [63:0] _current_y_5_T_7 = $signed(current_y_4) + $signed(_GEN_62); // @[Cordic_CR.scala 69:42]
  wire [63:0] _current_theta_5_T_5 = $signed(current_theta_4) - 64'sh1ca3794e5; // @[Cordic_CR.scala 70:50]
  wire [57:0] _current_x_6_T = current_y_5[63:6]; // @[Cordic_CR.scala 64:62]
  wire [63:0] _GEN_65 = {{6{_current_x_6_T[57]}},_current_x_6_T}; // @[Cordic_CR.scala 64:42]
  wire [63:0] _current_x_6_T_3 = $signed(current_x_5) + $signed(_GEN_65); // @[Cordic_CR.scala 64:42]
  wire [57:0] _current_y_6_T = current_x_5[63:6]; // @[Cordic_CR.scala 65:62]
  wire [63:0] _GEN_66 = {{6{_current_y_6_T[57]}},_current_y_6_T}; // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_y_6_T_3 = $signed(current_y_5) - $signed(_GEN_66); // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_theta_6_T_2 = $signed(current_theta_5) + 64'she52a1ab2; // @[Cordic_CR.scala 66:50]
  wire [63:0] _current_x_6_T_7 = $signed(current_x_5) - $signed(_GEN_65); // @[Cordic_CR.scala 68:42]
  wire [63:0] _current_y_6_T_7 = $signed(current_y_5) + $signed(_GEN_66); // @[Cordic_CR.scala 69:42]
  wire [63:0] _current_theta_6_T_5 = $signed(current_theta_5) - 64'she52a1ab2; // @[Cordic_CR.scala 70:50]
  wire [56:0] _current_x_7_T = current_y_6[63:7]; // @[Cordic_CR.scala 64:62]
  wire [63:0] _GEN_69 = {{7{_current_x_7_T[56]}},_current_x_7_T}; // @[Cordic_CR.scala 64:42]
  wire [63:0] _current_x_7_T_3 = $signed(current_x_6) + $signed(_GEN_69); // @[Cordic_CR.scala 64:42]
  wire [56:0] _current_y_7_T = current_x_6[63:7]; // @[Cordic_CR.scala 65:62]
  wire [63:0] _GEN_70 = {{7{_current_y_7_T[56]}},_current_y_7_T}; // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_y_7_T_3 = $signed(current_y_6) - $signed(_GEN_70); // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_theta_7_T_2 = $signed(current_theta_6) + 64'sh7296d7a1; // @[Cordic_CR.scala 66:50]
  wire [63:0] _current_x_7_T_7 = $signed(current_x_6) - $signed(_GEN_69); // @[Cordic_CR.scala 68:42]
  wire [63:0] _current_y_7_T_7 = $signed(current_y_6) + $signed(_GEN_70); // @[Cordic_CR.scala 69:42]
  wire [63:0] _current_theta_7_T_5 = $signed(current_theta_6) - 64'sh7296d7a1; // @[Cordic_CR.scala 70:50]
  wire [55:0] _current_x_8_T = current_y_7[63:8]; // @[Cordic_CR.scala 64:62]
  wire [63:0] _GEN_73 = {{8{_current_x_8_T[55]}},_current_x_8_T}; // @[Cordic_CR.scala 64:42]
  wire [63:0] _current_x_8_T_3 = $signed(current_x_7) + $signed(_GEN_73); // @[Cordic_CR.scala 64:42]
  wire [55:0] _current_y_8_T = current_x_7[63:8]; // @[Cordic_CR.scala 65:62]
  wire [63:0] _GEN_74 = {{8{_current_y_8_T[55]}},_current_y_8_T}; // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_y_8_T_3 = $signed(current_y_7) - $signed(_GEN_74); // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_theta_8_T_2 = $signed(current_theta_7) + 64'sh394ba51c; // @[Cordic_CR.scala 66:50]
  wire [63:0] _current_x_8_T_7 = $signed(current_x_7) - $signed(_GEN_73); // @[Cordic_CR.scala 68:42]
  wire [63:0] _current_y_8_T_7 = $signed(current_y_7) + $signed(_GEN_74); // @[Cordic_CR.scala 69:42]
  wire [63:0] _current_theta_8_T_5 = $signed(current_theta_7) - 64'sh394ba51c; // @[Cordic_CR.scala 70:50]
  wire [54:0] _current_x_9_T = current_y_8[63:9]; // @[Cordic_CR.scala 64:62]
  wire [63:0] _GEN_77 = {{9{_current_x_9_T[54]}},_current_x_9_T}; // @[Cordic_CR.scala 64:42]
  wire [63:0] _current_x_9_T_3 = $signed(current_x_8) + $signed(_GEN_77); // @[Cordic_CR.scala 64:42]
  wire [54:0] _current_y_9_T = current_x_8[63:9]; // @[Cordic_CR.scala 65:62]
  wire [63:0] _GEN_78 = {{9{_current_y_9_T[54]}},_current_y_9_T}; // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_y_9_T_3 = $signed(current_y_8) - $signed(_GEN_78); // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_theta_9_T_2 = $signed(current_theta_8) + 64'sh1ca5d9b7; // @[Cordic_CR.scala 66:50]
  wire [63:0] _current_x_9_T_7 = $signed(current_x_8) - $signed(_GEN_77); // @[Cordic_CR.scala 68:42]
  wire [63:0] _current_y_9_T_7 = $signed(current_y_8) + $signed(_GEN_78); // @[Cordic_CR.scala 69:42]
  wire [63:0] _current_theta_9_T_5 = $signed(current_theta_8) - 64'sh1ca5d9b7; // @[Cordic_CR.scala 70:50]
  wire [53:0] _current_x_10_T = current_y_9[63:10]; // @[Cordic_CR.scala 64:62]
  wire [63:0] _GEN_81 = {{10{_current_x_10_T[53]}},_current_x_10_T}; // @[Cordic_CR.scala 64:42]
  wire [63:0] _current_x_10_T_3 = $signed(current_x_9) + $signed(_GEN_81); // @[Cordic_CR.scala 64:42]
  wire [53:0] _current_y_10_T = current_x_9[63:10]; // @[Cordic_CR.scala 65:62]
  wire [63:0] _GEN_82 = {{10{_current_y_10_T[53]}},_current_y_10_T}; // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_y_10_T_3 = $signed(current_y_9) - $signed(_GEN_82); // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_theta_10_T_2 = $signed(current_theta_9) + 64'she52edc1; // @[Cordic_CR.scala 66:50]
  wire [63:0] _current_x_10_T_7 = $signed(current_x_9) - $signed(_GEN_81); // @[Cordic_CR.scala 68:42]
  wire [63:0] _current_y_10_T_7 = $signed(current_y_9) + $signed(_GEN_82); // @[Cordic_CR.scala 69:42]
  wire [63:0] _current_theta_10_T_5 = $signed(current_theta_9) - 64'she52edc1; // @[Cordic_CR.scala 70:50]
  wire [52:0] _current_x_11_T = current_y_10[63:11]; // @[Cordic_CR.scala 64:62]
  wire [63:0] _GEN_85 = {{11{_current_x_11_T[52]}},_current_x_11_T}; // @[Cordic_CR.scala 64:42]
  wire [63:0] _current_x_11_T_3 = $signed(current_x_10) + $signed(_GEN_85); // @[Cordic_CR.scala 64:42]
  wire [52:0] _current_y_11_T = current_x_10[63:11]; // @[Cordic_CR.scala 65:62]
  wire [63:0] _GEN_86 = {{11{_current_y_11_T[52]}},_current_y_11_T}; // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_y_11_T_3 = $signed(current_y_10) - $signed(_GEN_86); // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_theta_11_T_2 = $signed(current_theta_10) + 64'sh72976fd; // @[Cordic_CR.scala 66:50]
  wire [63:0] _current_x_11_T_7 = $signed(current_x_10) - $signed(_GEN_85); // @[Cordic_CR.scala 68:42]
  wire [63:0] _current_y_11_T_7 = $signed(current_y_10) + $signed(_GEN_86); // @[Cordic_CR.scala 69:42]
  wire [63:0] _current_theta_11_T_5 = $signed(current_theta_10) - 64'sh72976fd; // @[Cordic_CR.scala 70:50]
  wire [51:0] _current_x_12_T = current_y_11[63:12]; // @[Cordic_CR.scala 64:62]
  wire [63:0] _GEN_89 = {{12{_current_x_12_T[51]}},_current_x_12_T}; // @[Cordic_CR.scala 64:42]
  wire [63:0] _current_x_12_T_3 = $signed(current_x_11) + $signed(_GEN_89); // @[Cordic_CR.scala 64:42]
  wire [51:0] _current_y_12_T = current_x_11[63:12]; // @[Cordic_CR.scala 65:62]
  wire [63:0] _GEN_90 = {{12{_current_y_12_T[51]}},_current_y_12_T}; // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_y_12_T_3 = $signed(current_y_11) - $signed(_GEN_90); // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_theta_12_T_2 = $signed(current_theta_11) + 64'sh394bb82; // @[Cordic_CR.scala 66:50]
  wire [63:0] _current_x_12_T_7 = $signed(current_x_11) - $signed(_GEN_89); // @[Cordic_CR.scala 68:42]
  wire [63:0] _current_y_12_T_7 = $signed(current_y_11) + $signed(_GEN_90); // @[Cordic_CR.scala 69:42]
  wire [63:0] _current_theta_12_T_5 = $signed(current_theta_11) - 64'sh394bb82; // @[Cordic_CR.scala 70:50]
  wire [50:0] _current_x_13_T = current_y_12[63:13]; // @[Cordic_CR.scala 64:62]
  wire [63:0] _GEN_93 = {{13{_current_x_13_T[50]}},_current_x_13_T}; // @[Cordic_CR.scala 64:42]
  wire [63:0] _current_x_13_T_3 = $signed(current_x_12) + $signed(_GEN_93); // @[Cordic_CR.scala 64:42]
  wire [50:0] _current_y_13_T = current_x_12[63:13]; // @[Cordic_CR.scala 65:62]
  wire [63:0] _GEN_94 = {{13{_current_y_13_T[50]}},_current_y_13_T}; // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_y_13_T_3 = $signed(current_y_12) - $signed(_GEN_94); // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_theta_13_T_2 = $signed(current_theta_12) + 64'sh1ca5dc2; // @[Cordic_CR.scala 66:50]
  wire [63:0] _current_x_13_T_7 = $signed(current_x_12) - $signed(_GEN_93); // @[Cordic_CR.scala 68:42]
  wire [63:0] _current_y_13_T_7 = $signed(current_y_12) + $signed(_GEN_94); // @[Cordic_CR.scala 69:42]
  wire [63:0] _current_theta_13_T_5 = $signed(current_theta_12) - 64'sh1ca5dc2; // @[Cordic_CR.scala 70:50]
  wire [49:0] _current_x_14_T = current_y_13[63:14]; // @[Cordic_CR.scala 64:62]
  wire [63:0] _GEN_97 = {{14{_current_x_14_T[49]}},_current_x_14_T}; // @[Cordic_CR.scala 64:42]
  wire [63:0] _current_x_14_T_3 = $signed(current_x_13) + $signed(_GEN_97); // @[Cordic_CR.scala 64:42]
  wire [49:0] _current_y_14_T = current_x_13[63:14]; // @[Cordic_CR.scala 65:62]
  wire [63:0] _GEN_98 = {{14{_current_y_14_T[49]}},_current_y_14_T}; // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_y_14_T_3 = $signed(current_y_13) - $signed(_GEN_98); // @[Cordic_CR.scala 65:42]
  wire [63:0] _current_x_14_T_7 = $signed(current_x_13) - $signed(_GEN_97); // @[Cordic_CR.scala 68:42]
  wire [63:0] _current_y_14_T_7 = $signed(current_y_13) + $signed(_GEN_98); // @[Cordic_CR.scala 69:42]
  wire [127:0] _io_x_n_T = $signed(current_x_14) * 64'sh9b74eda8; // @[Cordic_CR.scala 80:43]
  wire [127:0] _io_y_n_T = $signed(current_y_14) * 64'sh9b74eda8; // @[Cordic_CR.scala 81:43]
  wire [95:0] _GEN_101 = _io_x_n_T[127:32]; // @[Cordic_CR.scala 80:10]
  wire [95:0] _GEN_103 = _io_y_n_T[127:32]; // @[Cordic_CR.scala 81:10]
  assign io_x_n = _GEN_101[63:0]; // @[Cordic_CR.scala 80:10]
  assign io_y_n = _GEN_103[63:0]; // @[Cordic_CR.scala 81:10]
  always @(posedge clock) begin
    if (reset) begin // @[Cordic_CR.scala 42:43]
      current_x_0 <= 64'sh0; // @[Cordic_CR.scala 42:43]
    end else if ($signed(io_theta) < 64'sh0) begin // @[Cordic_CR.scala 53:80]
      current_x_0 <= _current_x_0_T_2; // @[Cordic_CR.scala 54:22]
    end else begin
      current_x_0 <= _current_x_0_T_5; // @[Cordic_CR.scala 58:22]
    end
    if (reset) begin // @[Cordic_CR.scala 42:43]
      current_x_1 <= 64'sh0; // @[Cordic_CR.scala 42:43]
    end else if ($signed(current_theta_0) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_x_1 <= _current_x_1_T_3; // @[Cordic_CR.scala 64:22]
    end else begin
      current_x_1 <= _current_x_1_T_7; // @[Cordic_CR.scala 68:22]
    end
    if (reset) begin // @[Cordic_CR.scala 42:43]
      current_x_2 <= 64'sh0; // @[Cordic_CR.scala 42:43]
    end else if ($signed(current_theta_1) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_x_2 <= _current_x_2_T_3; // @[Cordic_CR.scala 64:22]
    end else begin
      current_x_2 <= _current_x_2_T_7; // @[Cordic_CR.scala 68:22]
    end
    if (reset) begin // @[Cordic_CR.scala 42:43]
      current_x_3 <= 64'sh0; // @[Cordic_CR.scala 42:43]
    end else if ($signed(current_theta_2) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_x_3 <= _current_x_3_T_3; // @[Cordic_CR.scala 64:22]
    end else begin
      current_x_3 <= _current_x_3_T_7; // @[Cordic_CR.scala 68:22]
    end
    if (reset) begin // @[Cordic_CR.scala 42:43]
      current_x_4 <= 64'sh0; // @[Cordic_CR.scala 42:43]
    end else if ($signed(current_theta_3) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_x_4 <= _current_x_4_T_3; // @[Cordic_CR.scala 64:22]
    end else begin
      current_x_4 <= _current_x_4_T_7; // @[Cordic_CR.scala 68:22]
    end
    if (reset) begin // @[Cordic_CR.scala 42:43]
      current_x_5 <= 64'sh0; // @[Cordic_CR.scala 42:43]
    end else if ($signed(current_theta_4) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_x_5 <= _current_x_5_T_3; // @[Cordic_CR.scala 64:22]
    end else begin
      current_x_5 <= _current_x_5_T_7; // @[Cordic_CR.scala 68:22]
    end
    if (reset) begin // @[Cordic_CR.scala 42:43]
      current_x_6 <= 64'sh0; // @[Cordic_CR.scala 42:43]
    end else if ($signed(current_theta_5) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_x_6 <= _current_x_6_T_3; // @[Cordic_CR.scala 64:22]
    end else begin
      current_x_6 <= _current_x_6_T_7; // @[Cordic_CR.scala 68:22]
    end
    if (reset) begin // @[Cordic_CR.scala 42:43]
      current_x_7 <= 64'sh0; // @[Cordic_CR.scala 42:43]
    end else if ($signed(current_theta_6) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_x_7 <= _current_x_7_T_3; // @[Cordic_CR.scala 64:22]
    end else begin
      current_x_7 <= _current_x_7_T_7; // @[Cordic_CR.scala 68:22]
    end
    if (reset) begin // @[Cordic_CR.scala 42:43]
      current_x_8 <= 64'sh0; // @[Cordic_CR.scala 42:43]
    end else if ($signed(current_theta_7) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_x_8 <= _current_x_8_T_3; // @[Cordic_CR.scala 64:22]
    end else begin
      current_x_8 <= _current_x_8_T_7; // @[Cordic_CR.scala 68:22]
    end
    if (reset) begin // @[Cordic_CR.scala 42:43]
      current_x_9 <= 64'sh0; // @[Cordic_CR.scala 42:43]
    end else if ($signed(current_theta_8) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_x_9 <= _current_x_9_T_3; // @[Cordic_CR.scala 64:22]
    end else begin
      current_x_9 <= _current_x_9_T_7; // @[Cordic_CR.scala 68:22]
    end
    if (reset) begin // @[Cordic_CR.scala 42:43]
      current_x_10 <= 64'sh0; // @[Cordic_CR.scala 42:43]
    end else if ($signed(current_theta_9) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_x_10 <= _current_x_10_T_3; // @[Cordic_CR.scala 64:22]
    end else begin
      current_x_10 <= _current_x_10_T_7; // @[Cordic_CR.scala 68:22]
    end
    if (reset) begin // @[Cordic_CR.scala 42:43]
      current_x_11 <= 64'sh0; // @[Cordic_CR.scala 42:43]
    end else if ($signed(current_theta_10) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_x_11 <= _current_x_11_T_3; // @[Cordic_CR.scala 64:22]
    end else begin
      current_x_11 <= _current_x_11_T_7; // @[Cordic_CR.scala 68:22]
    end
    if (reset) begin // @[Cordic_CR.scala 42:43]
      current_x_12 <= 64'sh0; // @[Cordic_CR.scala 42:43]
    end else if ($signed(current_theta_11) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_x_12 <= _current_x_12_T_3; // @[Cordic_CR.scala 64:22]
    end else begin
      current_x_12 <= _current_x_12_T_7; // @[Cordic_CR.scala 68:22]
    end
    if (reset) begin // @[Cordic_CR.scala 42:43]
      current_x_13 <= 64'sh0; // @[Cordic_CR.scala 42:43]
    end else if ($signed(current_theta_12) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_x_13 <= _current_x_13_T_3; // @[Cordic_CR.scala 64:22]
    end else begin
      current_x_13 <= _current_x_13_T_7; // @[Cordic_CR.scala 68:22]
    end
    if (reset) begin // @[Cordic_CR.scala 42:43]
      current_x_14 <= 64'sh0; // @[Cordic_CR.scala 42:43]
    end else if ($signed(current_theta_13) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_x_14 <= _current_x_14_T_3; // @[Cordic_CR.scala 64:22]
    end else begin
      current_x_14 <= _current_x_14_T_7; // @[Cordic_CR.scala 68:22]
    end
    if (reset) begin // @[Cordic_CR.scala 43:43]
      current_y_0 <= 64'sh0; // @[Cordic_CR.scala 43:43]
    end else if ($signed(io_theta) < 64'sh0) begin // @[Cordic_CR.scala 53:80]
      current_y_0 <= _current_y_0_T_5; // @[Cordic_CR.scala 55:22]
    end else begin
      current_y_0 <= _current_x_0_T_2; // @[Cordic_CR.scala 59:22]
    end
    if (reset) begin // @[Cordic_CR.scala 43:43]
      current_y_1 <= 64'sh0; // @[Cordic_CR.scala 43:43]
    end else if ($signed(current_theta_0) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_y_1 <= _current_y_1_T_3; // @[Cordic_CR.scala 65:22]
    end else begin
      current_y_1 <= _current_y_1_T_7; // @[Cordic_CR.scala 69:22]
    end
    if (reset) begin // @[Cordic_CR.scala 43:43]
      current_y_2 <= 64'sh0; // @[Cordic_CR.scala 43:43]
    end else if ($signed(current_theta_1) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_y_2 <= _current_y_2_T_3; // @[Cordic_CR.scala 65:22]
    end else begin
      current_y_2 <= _current_y_2_T_7; // @[Cordic_CR.scala 69:22]
    end
    if (reset) begin // @[Cordic_CR.scala 43:43]
      current_y_3 <= 64'sh0; // @[Cordic_CR.scala 43:43]
    end else if ($signed(current_theta_2) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_y_3 <= _current_y_3_T_3; // @[Cordic_CR.scala 65:22]
    end else begin
      current_y_3 <= _current_y_3_T_7; // @[Cordic_CR.scala 69:22]
    end
    if (reset) begin // @[Cordic_CR.scala 43:43]
      current_y_4 <= 64'sh0; // @[Cordic_CR.scala 43:43]
    end else if ($signed(current_theta_3) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_y_4 <= _current_y_4_T_3; // @[Cordic_CR.scala 65:22]
    end else begin
      current_y_4 <= _current_y_4_T_7; // @[Cordic_CR.scala 69:22]
    end
    if (reset) begin // @[Cordic_CR.scala 43:43]
      current_y_5 <= 64'sh0; // @[Cordic_CR.scala 43:43]
    end else if ($signed(current_theta_4) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_y_5 <= _current_y_5_T_3; // @[Cordic_CR.scala 65:22]
    end else begin
      current_y_5 <= _current_y_5_T_7; // @[Cordic_CR.scala 69:22]
    end
    if (reset) begin // @[Cordic_CR.scala 43:43]
      current_y_6 <= 64'sh0; // @[Cordic_CR.scala 43:43]
    end else if ($signed(current_theta_5) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_y_6 <= _current_y_6_T_3; // @[Cordic_CR.scala 65:22]
    end else begin
      current_y_6 <= _current_y_6_T_7; // @[Cordic_CR.scala 69:22]
    end
    if (reset) begin // @[Cordic_CR.scala 43:43]
      current_y_7 <= 64'sh0; // @[Cordic_CR.scala 43:43]
    end else if ($signed(current_theta_6) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_y_7 <= _current_y_7_T_3; // @[Cordic_CR.scala 65:22]
    end else begin
      current_y_7 <= _current_y_7_T_7; // @[Cordic_CR.scala 69:22]
    end
    if (reset) begin // @[Cordic_CR.scala 43:43]
      current_y_8 <= 64'sh0; // @[Cordic_CR.scala 43:43]
    end else if ($signed(current_theta_7) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_y_8 <= _current_y_8_T_3; // @[Cordic_CR.scala 65:22]
    end else begin
      current_y_8 <= _current_y_8_T_7; // @[Cordic_CR.scala 69:22]
    end
    if (reset) begin // @[Cordic_CR.scala 43:43]
      current_y_9 <= 64'sh0; // @[Cordic_CR.scala 43:43]
    end else if ($signed(current_theta_8) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_y_9 <= _current_y_9_T_3; // @[Cordic_CR.scala 65:22]
    end else begin
      current_y_9 <= _current_y_9_T_7; // @[Cordic_CR.scala 69:22]
    end
    if (reset) begin // @[Cordic_CR.scala 43:43]
      current_y_10 <= 64'sh0; // @[Cordic_CR.scala 43:43]
    end else if ($signed(current_theta_9) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_y_10 <= _current_y_10_T_3; // @[Cordic_CR.scala 65:22]
    end else begin
      current_y_10 <= _current_y_10_T_7; // @[Cordic_CR.scala 69:22]
    end
    if (reset) begin // @[Cordic_CR.scala 43:43]
      current_y_11 <= 64'sh0; // @[Cordic_CR.scala 43:43]
    end else if ($signed(current_theta_10) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_y_11 <= _current_y_11_T_3; // @[Cordic_CR.scala 65:22]
    end else begin
      current_y_11 <= _current_y_11_T_7; // @[Cordic_CR.scala 69:22]
    end
    if (reset) begin // @[Cordic_CR.scala 43:43]
      current_y_12 <= 64'sh0; // @[Cordic_CR.scala 43:43]
    end else if ($signed(current_theta_11) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_y_12 <= _current_y_12_T_3; // @[Cordic_CR.scala 65:22]
    end else begin
      current_y_12 <= _current_y_12_T_7; // @[Cordic_CR.scala 69:22]
    end
    if (reset) begin // @[Cordic_CR.scala 43:43]
      current_y_13 <= 64'sh0; // @[Cordic_CR.scala 43:43]
    end else if ($signed(current_theta_12) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_y_13 <= _current_y_13_T_3; // @[Cordic_CR.scala 65:22]
    end else begin
      current_y_13 <= _current_y_13_T_7; // @[Cordic_CR.scala 69:22]
    end
    if (reset) begin // @[Cordic_CR.scala 43:43]
      current_y_14 <= 64'sh0; // @[Cordic_CR.scala 43:43]
    end else if ($signed(current_theta_13) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_y_14 <= _current_y_14_T_3; // @[Cordic_CR.scala 65:22]
    end else begin
      current_y_14 <= _current_y_14_T_7; // @[Cordic_CR.scala 69:22]
    end
    if (reset) begin // @[Cordic_CR.scala 44:47]
      current_theta_0 <= 64'sh0; // @[Cordic_CR.scala 44:47]
    end else if ($signed(io_theta) < 64'sh0) begin // @[Cordic_CR.scala 53:80]
      current_theta_0 <= _current_theta_0_T_2; // @[Cordic_CR.scala 56:26]
    end else begin
      current_theta_0 <= _current_theta_0_T_5; // @[Cordic_CR.scala 60:26]
    end
    if (reset) begin // @[Cordic_CR.scala 44:47]
      current_theta_1 <= 64'sh0; // @[Cordic_CR.scala 44:47]
    end else if ($signed(current_theta_0) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_theta_1 <= _current_theta_1_T_2; // @[Cordic_CR.scala 66:26]
    end else begin
      current_theta_1 <= _current_theta_1_T_5; // @[Cordic_CR.scala 70:26]
    end
    if (reset) begin // @[Cordic_CR.scala 44:47]
      current_theta_2 <= 64'sh0; // @[Cordic_CR.scala 44:47]
    end else if ($signed(current_theta_1) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_theta_2 <= _current_theta_2_T_2; // @[Cordic_CR.scala 66:26]
    end else begin
      current_theta_2 <= _current_theta_2_T_5; // @[Cordic_CR.scala 70:26]
    end
    if (reset) begin // @[Cordic_CR.scala 44:47]
      current_theta_3 <= 64'sh0; // @[Cordic_CR.scala 44:47]
    end else if ($signed(current_theta_2) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_theta_3 <= _current_theta_3_T_2; // @[Cordic_CR.scala 66:26]
    end else begin
      current_theta_3 <= _current_theta_3_T_5; // @[Cordic_CR.scala 70:26]
    end
    if (reset) begin // @[Cordic_CR.scala 44:47]
      current_theta_4 <= 64'sh0; // @[Cordic_CR.scala 44:47]
    end else if ($signed(current_theta_3) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_theta_4 <= _current_theta_4_T_2; // @[Cordic_CR.scala 66:26]
    end else begin
      current_theta_4 <= _current_theta_4_T_5; // @[Cordic_CR.scala 70:26]
    end
    if (reset) begin // @[Cordic_CR.scala 44:47]
      current_theta_5 <= 64'sh0; // @[Cordic_CR.scala 44:47]
    end else if ($signed(current_theta_4) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_theta_5 <= _current_theta_5_T_2; // @[Cordic_CR.scala 66:26]
    end else begin
      current_theta_5 <= _current_theta_5_T_5; // @[Cordic_CR.scala 70:26]
    end
    if (reset) begin // @[Cordic_CR.scala 44:47]
      current_theta_6 <= 64'sh0; // @[Cordic_CR.scala 44:47]
    end else if ($signed(current_theta_5) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_theta_6 <= _current_theta_6_T_2; // @[Cordic_CR.scala 66:26]
    end else begin
      current_theta_6 <= _current_theta_6_T_5; // @[Cordic_CR.scala 70:26]
    end
    if (reset) begin // @[Cordic_CR.scala 44:47]
      current_theta_7 <= 64'sh0; // @[Cordic_CR.scala 44:47]
    end else if ($signed(current_theta_6) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_theta_7 <= _current_theta_7_T_2; // @[Cordic_CR.scala 66:26]
    end else begin
      current_theta_7 <= _current_theta_7_T_5; // @[Cordic_CR.scala 70:26]
    end
    if (reset) begin // @[Cordic_CR.scala 44:47]
      current_theta_8 <= 64'sh0; // @[Cordic_CR.scala 44:47]
    end else if ($signed(current_theta_7) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_theta_8 <= _current_theta_8_T_2; // @[Cordic_CR.scala 66:26]
    end else begin
      current_theta_8 <= _current_theta_8_T_5; // @[Cordic_CR.scala 70:26]
    end
    if (reset) begin // @[Cordic_CR.scala 44:47]
      current_theta_9 <= 64'sh0; // @[Cordic_CR.scala 44:47]
    end else if ($signed(current_theta_8) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_theta_9 <= _current_theta_9_T_2; // @[Cordic_CR.scala 66:26]
    end else begin
      current_theta_9 <= _current_theta_9_T_5; // @[Cordic_CR.scala 70:26]
    end
    if (reset) begin // @[Cordic_CR.scala 44:47]
      current_theta_10 <= 64'sh0; // @[Cordic_CR.scala 44:47]
    end else if ($signed(current_theta_9) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_theta_10 <= _current_theta_10_T_2; // @[Cordic_CR.scala 66:26]
    end else begin
      current_theta_10 <= _current_theta_10_T_5; // @[Cordic_CR.scala 70:26]
    end
    if (reset) begin // @[Cordic_CR.scala 44:47]
      current_theta_11 <= 64'sh0; // @[Cordic_CR.scala 44:47]
    end else if ($signed(current_theta_10) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_theta_11 <= _current_theta_11_T_2; // @[Cordic_CR.scala 66:26]
    end else begin
      current_theta_11 <= _current_theta_11_T_5; // @[Cordic_CR.scala 70:26]
    end
    if (reset) begin // @[Cordic_CR.scala 44:47]
      current_theta_12 <= 64'sh0; // @[Cordic_CR.scala 44:47]
    end else if ($signed(current_theta_11) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_theta_12 <= _current_theta_12_T_2; // @[Cordic_CR.scala 66:26]
    end else begin
      current_theta_12 <= _current_theta_12_T_5; // @[Cordic_CR.scala 70:26]
    end
    if (reset) begin // @[Cordic_CR.scala 44:47]
      current_theta_13 <= 64'sh0; // @[Cordic_CR.scala 44:47]
    end else if ($signed(current_theta_12) < 64'sh0) begin // @[Cordic_CR.scala 63:92]
      current_theta_13 <= _current_theta_13_T_2; // @[Cordic_CR.scala 66:26]
    end else begin
      current_theta_13 <= _current_theta_13_T_5; // @[Cordic_CR.scala 70:26]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  current_x_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  current_x_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  current_x_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  current_x_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  current_x_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  current_x_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  current_x_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  current_x_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  current_x_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  current_x_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  current_x_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  current_x_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  current_x_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  current_x_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  current_x_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  current_y_0 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  current_y_1 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  current_y_2 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  current_y_3 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  current_y_4 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  current_y_5 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  current_y_6 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  current_y_7 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  current_y_8 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  current_y_9 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  current_y_10 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  current_y_11 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  current_y_12 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  current_y_13 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  current_y_14 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  current_theta_0 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  current_theta_1 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  current_theta_2 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  current_theta_3 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  current_theta_4 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  current_theta_5 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  current_theta_6 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  current_theta_7 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  current_theta_8 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  current_theta_9 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  current_theta_10 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  current_theta_11 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  current_theta_12 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  current_theta_13 = _RAND_43[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cordic_sin_cos(
  input         clock,
  input         reset,
  input  [63:0] io_theta,
  output [63:0] io_sin,
  output [63:0] io_cos
);
  wire  cordic_unit_clock; // @[Cordic_CR.scala 145:45]
  wire  cordic_unit_reset; // @[Cordic_CR.scala 145:45]
  wire [63:0] cordic_unit_io_x; // @[Cordic_CR.scala 145:45]
  wire [63:0] cordic_unit_io_y; // @[Cordic_CR.scala 145:45]
  wire [63:0] cordic_unit_io_theta; // @[Cordic_CR.scala 145:45]
  wire [63:0] cordic_unit_io_x_n; // @[Cordic_CR.scala 145:45]
  wire [63:0] cordic_unit_io_y_n; // @[Cordic_CR.scala 145:45]
  wire [63:0] _temp_theta_T_2 = $signed(io_theta) - 64'sh16800000000; // @[Cordic_CR.scala 123:28]
  wire [63:0] _temp_theta_T_5 = $signed(io_theta) + 64'sh16800000000; // @[Cordic_CR.scala 125:28]
  wire [63:0] _GEN_0 = $signed(io_theta) < -64'shb400000000 ? $signed(_temp_theta_T_5) : $signed(io_theta); // @[Cordic_CR.scala 124:83 125:16 127:16]
  wire [63:0] temp_theta = $signed(io_theta) > 64'shb400000000 ? $signed(_temp_theta_T_2) : $signed(_GEN_0); // @[Cordic_CR.scala 122:76 123:16]
  wire  _T_2 = $signed(temp_theta) > 64'sh5a00000000; // @[Cordic_CR.scala 133:19]
  wire [63:0] _real_theta_T_2 = 64'shb400000000 - $signed(temp_theta); // @[Cordic_CR.scala 136:75]
  wire [63:0] _real_theta_T_5 = -64'shb400000000 - $signed(temp_theta); // @[Cordic_CR.scala 139:76]
  wire  _GEN_2 = $signed(temp_theta) < -64'sh5a00000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 137:84 138:15 141:15]
  wire [63:0] _GEN_3 = $signed(temp_theta) < -64'sh5a00000000 ? $signed(_real_theta_T_5) : $signed(temp_theta); // @[Cordic_CR.scala 137:84 139:16 142:16]
  wire  sigma_cos = _T_2 ? 1'h0 : _GEN_2; // @[Cordic_CR.scala 134:5 135:15]
  wire [63:0] _io_cos_T_2 = 64'sh0 - $signed(cordic_unit_io_x_n); // @[Cordic_CR.scala 153:15]
  CORDIC_CR_ORIGIN cordic_unit ( // @[Cordic_CR.scala 145:45]
    .clock(cordic_unit_clock),
    .reset(cordic_unit_reset),
    .io_x(cordic_unit_io_x),
    .io_y(cordic_unit_io_y),
    .io_theta(cordic_unit_io_theta),
    .io_x_n(cordic_unit_io_x_n),
    .io_y_n(cordic_unit_io_y_n)
  );
  assign io_sin = cordic_unit_io_y_n; // @[Cordic_CR.scala 149:10]
  assign io_cos = sigma_cos ? $signed(cordic_unit_io_x_n) : $signed(_io_cos_T_2); // @[Cordic_CR.scala 150:19 151:12 153:12]
  assign cordic_unit_clock = clock;
  assign cordic_unit_reset = reset;
  assign cordic_unit_io_x = 64'sh100000000; // @[Cordic_CR.scala 146:20]
  assign cordic_unit_io_y = 64'sh0; // @[Cordic_CR.scala 147:20]
  assign cordic_unit_io_theta = _T_2 ? $signed(_real_theta_T_2) : $signed(_GEN_3); // @[Cordic_CR.scala 134:5 136:16]
endmodule
module shift_2_range(
  input  [63:0] io_x,
  output [63:0] io_out,
  output [5:0]  io_cnt,
  output        io_flag
);
  wire [63:0] _temp_x_T_2 = 64'sh0 - $signed(io_x); // @[Cordic_LV.scala 77:15]
  wire [63:0] temp_x = $signed(io_x) < 64'sh0 ? $signed(_temp_x_T_2) : $signed(io_x); // @[Cordic_LV.scala 76:72 77:12 80:12]
  wire  _T_1 = $signed(temp_x) < 64'sh80000000; // @[Cordic_LV.scala 84:15]
  wire  index__0 = _T_1 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [64:0] _T_4 = {$signed(temp_x), 1'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__1 = $signed(_T_4) < 65'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [65:0] _T_6 = {$signed(temp_x), 2'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__2 = $signed(_T_6) < 66'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [66:0] _T_8 = {$signed(temp_x), 3'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__3 = $signed(_T_8) < 67'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [67:0] _T_10 = {$signed(temp_x), 4'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__4 = $signed(_T_10) < 68'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [68:0] _T_12 = {$signed(temp_x), 5'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__5 = $signed(_T_12) < 69'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [69:0] _T_14 = {$signed(temp_x), 6'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__6 = $signed(_T_14) < 70'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [70:0] _T_16 = {$signed(temp_x), 7'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__7 = $signed(_T_16) < 71'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [71:0] _T_18 = {$signed(temp_x), 8'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__8 = $signed(_T_18) < 72'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [72:0] _T_20 = {$signed(temp_x), 9'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__9 = $signed(_T_20) < 73'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [73:0] _T_22 = {$signed(temp_x), 10'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__10 = $signed(_T_22) < 74'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [74:0] _T_24 = {$signed(temp_x), 11'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__11 = $signed(_T_24) < 75'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [75:0] _T_26 = {$signed(temp_x), 12'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__12 = $signed(_T_26) < 76'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [76:0] _T_28 = {$signed(temp_x), 13'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__13 = $signed(_T_28) < 77'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [77:0] _T_30 = {$signed(temp_x), 14'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__14 = $signed(_T_30) < 78'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [78:0] _T_32 = {$signed(temp_x), 15'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__15 = $signed(_T_32) < 79'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [79:0] _T_34 = {$signed(temp_x), 16'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__16 = $signed(_T_34) < 80'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [80:0] _T_36 = {$signed(temp_x), 17'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__17 = $signed(_T_36) < 81'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [81:0] _T_38 = {$signed(temp_x), 18'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__18 = $signed(_T_38) < 82'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [82:0] _T_40 = {$signed(temp_x), 19'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__19 = $signed(_T_40) < 83'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [83:0] _T_42 = {$signed(temp_x), 20'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__20 = $signed(_T_42) < 84'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [84:0] _T_44 = {$signed(temp_x), 21'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__21 = $signed(_T_44) < 85'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [85:0] _T_46 = {$signed(temp_x), 22'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__22 = $signed(_T_46) < 86'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [86:0] _T_48 = {$signed(temp_x), 23'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__23 = $signed(_T_48) < 87'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [87:0] _T_50 = {$signed(temp_x), 24'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__24 = $signed(_T_50) < 88'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [88:0] _T_52 = {$signed(temp_x), 25'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__25 = $signed(_T_52) < 89'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [89:0] _T_54 = {$signed(temp_x), 26'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__26 = $signed(_T_54) < 90'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [90:0] _T_56 = {$signed(temp_x), 27'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__27 = $signed(_T_56) < 91'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [91:0] _T_58 = {$signed(temp_x), 28'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__28 = $signed(_T_58) < 92'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [92:0] _T_60 = {$signed(temp_x), 29'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__29 = $signed(_T_60) < 93'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [93:0] _T_62 = {$signed(temp_x), 30'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__30 = $signed(_T_62) < 94'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [94:0] _T_64 = {$signed(temp_x), 31'h0}; // @[Cordic_LV.scala 88:20]
  wire  index__31 = $signed(_T_64) < 95'sh80000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 88:85 89:18 91:18]
  wire [7:0] temp_cnt_lo_lo = {index__7,index__6,index__5,index__4,index__3,index__2,index__1,index__0}; // @[Cordic_LV.scala 95:48]
  wire [15:0] temp_cnt_lo = {index__15,index__14,index__13,index__12,index__11,index__10,index__9,index__8,
    temp_cnt_lo_lo}; // @[Cordic_LV.scala 95:48]
  wire [7:0] temp_cnt_hi_lo = {index__23,index__22,index__21,index__20,index__19,index__18,index__17,index__16}; // @[Cordic_LV.scala 95:48]
  wire [31:0] _temp_cnt_T = {index__31,index__30,index__29,index__28,index__27,index__26,index__25,index__24,
    temp_cnt_hi_lo,temp_cnt_lo}; // @[Cordic_LV.scala 95:48]
  wire [4:0] _temp_cnt_T_33 = _temp_cnt_T[30] ? 5'h1e : 5'h1f; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_34 = _temp_cnt_T[29] ? 5'h1d : _temp_cnt_T_33; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_35 = _temp_cnt_T[28] ? 5'h1c : _temp_cnt_T_34; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_36 = _temp_cnt_T[27] ? 5'h1b : _temp_cnt_T_35; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_37 = _temp_cnt_T[26] ? 5'h1a : _temp_cnt_T_36; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_38 = _temp_cnt_T[25] ? 5'h19 : _temp_cnt_T_37; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_39 = _temp_cnt_T[24] ? 5'h18 : _temp_cnt_T_38; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_40 = _temp_cnt_T[23] ? 5'h17 : _temp_cnt_T_39; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_41 = _temp_cnt_T[22] ? 5'h16 : _temp_cnt_T_40; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_42 = _temp_cnt_T[21] ? 5'h15 : _temp_cnt_T_41; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_43 = _temp_cnt_T[20] ? 5'h14 : _temp_cnt_T_42; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_44 = _temp_cnt_T[19] ? 5'h13 : _temp_cnt_T_43; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_45 = _temp_cnt_T[18] ? 5'h12 : _temp_cnt_T_44; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_46 = _temp_cnt_T[17] ? 5'h11 : _temp_cnt_T_45; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_47 = _temp_cnt_T[16] ? 5'h10 : _temp_cnt_T_46; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_48 = _temp_cnt_T[15] ? 5'hf : _temp_cnt_T_47; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_49 = _temp_cnt_T[14] ? 5'he : _temp_cnt_T_48; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_50 = _temp_cnt_T[13] ? 5'hd : _temp_cnt_T_49; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_51 = _temp_cnt_T[12] ? 5'hc : _temp_cnt_T_50; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_52 = _temp_cnt_T[11] ? 5'hb : _temp_cnt_T_51; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_53 = _temp_cnt_T[10] ? 5'ha : _temp_cnt_T_52; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_54 = _temp_cnt_T[9] ? 5'h9 : _temp_cnt_T_53; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_55 = _temp_cnt_T[8] ? 5'h8 : _temp_cnt_T_54; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_56 = _temp_cnt_T[7] ? 5'h7 : _temp_cnt_T_55; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_57 = _temp_cnt_T[6] ? 5'h6 : _temp_cnt_T_56; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_58 = _temp_cnt_T[5] ? 5'h5 : _temp_cnt_T_57; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_59 = _temp_cnt_T[4] ? 5'h4 : _temp_cnt_T_58; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_60 = _temp_cnt_T[3] ? 5'h3 : _temp_cnt_T_59; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_61 = _temp_cnt_T[2] ? 5'h2 : _temp_cnt_T_60; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_62 = _temp_cnt_T[1] ? 5'h1 : _temp_cnt_T_61; // @[Mux.scala 47:70]
  wire [4:0] temp_cnt = _temp_cnt_T[0] ? 5'h0 : _temp_cnt_T_62; // @[Mux.scala 47:70]
  wire [4:0] _io_cnt_T = _temp_cnt_T[0] ? 5'h0 : _temp_cnt_T_62; // @[Cordic_LV.scala 96:30]
  wire [94:0] _GEN_0 = {{31{temp_x[63]}},temp_x}; // @[Cordic_LV.scala 97:23]
  wire [94:0] _io_out_T = $signed(_GEN_0) << temp_cnt; // @[Cordic_LV.scala 97:23]
  wire  _T_66 = $signed(temp_x) > 64'sh100000000; // @[Cordic_LV.scala 98:21]
  wire  index_1_0 = _T_66 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [62:0] _T_69 = temp_x[63:1]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_102 = {{1{_T_69[62]}},_T_69}; // @[Cordic_LV.scala 102:26]
  wire  index_1_1 = $signed(_GEN_102) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [61:0] _T_71 = temp_x[63:2]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_103 = {{2{_T_71[61]}},_T_71}; // @[Cordic_LV.scala 102:26]
  wire  index_1_2 = $signed(_GEN_103) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [60:0] _T_73 = temp_x[63:3]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_104 = {{3{_T_73[60]}},_T_73}; // @[Cordic_LV.scala 102:26]
  wire  index_1_3 = $signed(_GEN_104) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [59:0] _T_75 = temp_x[63:4]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_105 = {{4{_T_75[59]}},_T_75}; // @[Cordic_LV.scala 102:26]
  wire  index_1_4 = $signed(_GEN_105) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [58:0] _T_77 = temp_x[63:5]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_106 = {{5{_T_77[58]}},_T_77}; // @[Cordic_LV.scala 102:26]
  wire  index_1_5 = $signed(_GEN_106) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [57:0] _T_79 = temp_x[63:6]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_107 = {{6{_T_79[57]}},_T_79}; // @[Cordic_LV.scala 102:26]
  wire  index_1_6 = $signed(_GEN_107) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [56:0] _T_81 = temp_x[63:7]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_108 = {{7{_T_81[56]}},_T_81}; // @[Cordic_LV.scala 102:26]
  wire  index_1_7 = $signed(_GEN_108) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [55:0] _T_83 = temp_x[63:8]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_109 = {{8{_T_83[55]}},_T_83}; // @[Cordic_LV.scala 102:26]
  wire  index_1_8 = $signed(_GEN_109) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [54:0] _T_85 = temp_x[63:9]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_110 = {{9{_T_85[54]}},_T_85}; // @[Cordic_LV.scala 102:26]
  wire  index_1_9 = $signed(_GEN_110) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [53:0] _T_87 = temp_x[63:10]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_111 = {{10{_T_87[53]}},_T_87}; // @[Cordic_LV.scala 102:26]
  wire  index_1_10 = $signed(_GEN_111) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [52:0] _T_89 = temp_x[63:11]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_112 = {{11{_T_89[52]}},_T_89}; // @[Cordic_LV.scala 102:26]
  wire  index_1_11 = $signed(_GEN_112) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [51:0] _T_91 = temp_x[63:12]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_113 = {{12{_T_91[51]}},_T_91}; // @[Cordic_LV.scala 102:26]
  wire  index_1_12 = $signed(_GEN_113) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [50:0] _T_93 = temp_x[63:13]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_114 = {{13{_T_93[50]}},_T_93}; // @[Cordic_LV.scala 102:26]
  wire  index_1_13 = $signed(_GEN_114) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [49:0] _T_95 = temp_x[63:14]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_115 = {{14{_T_95[49]}},_T_95}; // @[Cordic_LV.scala 102:26]
  wire  index_1_14 = $signed(_GEN_115) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [48:0] _T_97 = temp_x[63:15]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_116 = {{15{_T_97[48]}},_T_97}; // @[Cordic_LV.scala 102:26]
  wire  index_1_15 = $signed(_GEN_116) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [47:0] _T_99 = temp_x[63:16]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_117 = {{16{_T_99[47]}},_T_99}; // @[Cordic_LV.scala 102:26]
  wire  index_1_16 = $signed(_GEN_117) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [46:0] _T_101 = temp_x[63:17]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_118 = {{17{_T_101[46]}},_T_101}; // @[Cordic_LV.scala 102:26]
  wire  index_1_17 = $signed(_GEN_118) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [45:0] _T_103 = temp_x[63:18]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_119 = {{18{_T_103[45]}},_T_103}; // @[Cordic_LV.scala 102:26]
  wire  index_1_18 = $signed(_GEN_119) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [44:0] _T_105 = temp_x[63:19]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_120 = {{19{_T_105[44]}},_T_105}; // @[Cordic_LV.scala 102:26]
  wire  index_1_19 = $signed(_GEN_120) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [43:0] _T_107 = temp_x[63:20]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_121 = {{20{_T_107[43]}},_T_107}; // @[Cordic_LV.scala 102:26]
  wire  index_1_20 = $signed(_GEN_121) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [42:0] _T_109 = temp_x[63:21]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_122 = {{21{_T_109[42]}},_T_109}; // @[Cordic_LV.scala 102:26]
  wire  index_1_21 = $signed(_GEN_122) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [41:0] _T_111 = temp_x[63:22]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_123 = {{22{_T_111[41]}},_T_111}; // @[Cordic_LV.scala 102:26]
  wire  index_1_22 = $signed(_GEN_123) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [40:0] _T_113 = temp_x[63:23]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_124 = {{23{_T_113[40]}},_T_113}; // @[Cordic_LV.scala 102:26]
  wire  index_1_23 = $signed(_GEN_124) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [39:0] _T_115 = temp_x[63:24]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_125 = {{24{_T_115[39]}},_T_115}; // @[Cordic_LV.scala 102:26]
  wire  index_1_24 = $signed(_GEN_125) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [38:0] _T_117 = temp_x[63:25]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_126 = {{25{_T_117[38]}},_T_117}; // @[Cordic_LV.scala 102:26]
  wire  index_1_25 = $signed(_GEN_126) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [37:0] _T_119 = temp_x[63:26]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_127 = {{26{_T_119[37]}},_T_119}; // @[Cordic_LV.scala 102:26]
  wire  index_1_26 = $signed(_GEN_127) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [36:0] _T_121 = temp_x[63:27]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_128 = {{27{_T_121[36]}},_T_121}; // @[Cordic_LV.scala 102:26]
  wire  index_1_27 = $signed(_GEN_128) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [35:0] _T_123 = temp_x[63:28]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_129 = {{28{_T_123[35]}},_T_123}; // @[Cordic_LV.scala 102:26]
  wire  index_1_28 = $signed(_GEN_129) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [34:0] _T_125 = temp_x[63:29]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_130 = {{29{_T_125[34]}},_T_125}; // @[Cordic_LV.scala 102:26]
  wire  index_1_29 = $signed(_GEN_130) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [33:0] _T_127 = temp_x[63:30]; // @[Cordic_LV.scala 102:20]
  wire [63:0] _GEN_131 = {{30{_T_127[33]}},_T_127}; // @[Cordic_LV.scala 102:26]
  wire  index_1_30 = $signed(_GEN_131) > 64'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 102:83 103:18 105:18]
  wire [7:0] temp_cnt_lo_lo_lo_1 = {index_1_7,index_1_6,index_1_5,index_1_4,index_1_3,index_1_2,index_1_1,index_1_0}; // @[Cordic_LV.scala 109:48]
  wire [15:0] temp_cnt_lo_lo_1 = {index_1_15,index_1_14,index_1_13,index_1_12,index_1_11,index_1_10,index_1_9,index_1_8,
    temp_cnt_lo_lo_lo_1}; // @[Cordic_LV.scala 109:48]
  wire [7:0] temp_cnt_lo_hi_lo_1 = {index_1_23,index_1_22,index_1_21,index_1_20,index_1_19,index_1_18,index_1_17,
    index_1_16}; // @[Cordic_LV.scala 109:48]
  wire [31:0] temp_cnt_lo_1 = {1'h1,index_1_30,index_1_29,index_1_28,index_1_27,index_1_26,index_1_25,index_1_24,
    temp_cnt_lo_hi_lo_1,temp_cnt_lo_lo_1}; // @[Cordic_LV.scala 109:48]
  wire [63:0] _temp_cnt_T_63 = {32'hffffffff,temp_cnt_lo_1}; // @[Cordic_LV.scala 109:48]
  wire [5:0] _temp_cnt_T_128 = _temp_cnt_T_63[62] ? 6'h3e : 6'h3f; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_129 = _temp_cnt_T_63[61] ? 6'h3d : _temp_cnt_T_128; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_130 = _temp_cnt_T_63[60] ? 6'h3c : _temp_cnt_T_129; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_131 = _temp_cnt_T_63[59] ? 6'h3b : _temp_cnt_T_130; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_132 = _temp_cnt_T_63[58] ? 6'h3a : _temp_cnt_T_131; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_133 = _temp_cnt_T_63[57] ? 6'h39 : _temp_cnt_T_132; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_134 = _temp_cnt_T_63[56] ? 6'h38 : _temp_cnt_T_133; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_135 = _temp_cnt_T_63[55] ? 6'h37 : _temp_cnt_T_134; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_136 = _temp_cnt_T_63[54] ? 6'h36 : _temp_cnt_T_135; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_137 = _temp_cnt_T_63[53] ? 6'h35 : _temp_cnt_T_136; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_138 = _temp_cnt_T_63[52] ? 6'h34 : _temp_cnt_T_137; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_139 = _temp_cnt_T_63[51] ? 6'h33 : _temp_cnt_T_138; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_140 = _temp_cnt_T_63[50] ? 6'h32 : _temp_cnt_T_139; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_141 = _temp_cnt_T_63[49] ? 6'h31 : _temp_cnt_T_140; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_142 = _temp_cnt_T_63[48] ? 6'h30 : _temp_cnt_T_141; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_143 = _temp_cnt_T_63[47] ? 6'h2f : _temp_cnt_T_142; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_144 = _temp_cnt_T_63[46] ? 6'h2e : _temp_cnt_T_143; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_145 = _temp_cnt_T_63[45] ? 6'h2d : _temp_cnt_T_144; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_146 = _temp_cnt_T_63[44] ? 6'h2c : _temp_cnt_T_145; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_147 = _temp_cnt_T_63[43] ? 6'h2b : _temp_cnt_T_146; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_148 = _temp_cnt_T_63[42] ? 6'h2a : _temp_cnt_T_147; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_149 = _temp_cnt_T_63[41] ? 6'h29 : _temp_cnt_T_148; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_150 = _temp_cnt_T_63[40] ? 6'h28 : _temp_cnt_T_149; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_151 = _temp_cnt_T_63[39] ? 6'h27 : _temp_cnt_T_150; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_152 = _temp_cnt_T_63[38] ? 6'h26 : _temp_cnt_T_151; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_153 = _temp_cnt_T_63[37] ? 6'h25 : _temp_cnt_T_152; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_154 = _temp_cnt_T_63[36] ? 6'h24 : _temp_cnt_T_153; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_155 = _temp_cnt_T_63[35] ? 6'h23 : _temp_cnt_T_154; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_156 = _temp_cnt_T_63[34] ? 6'h22 : _temp_cnt_T_155; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_157 = _temp_cnt_T_63[33] ? 6'h21 : _temp_cnt_T_156; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_158 = _temp_cnt_T_63[32] ? 6'h20 : _temp_cnt_T_157; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_159 = _temp_cnt_T_63[31] ? 6'h1f : _temp_cnt_T_158; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_160 = _temp_cnt_T_63[30] ? 6'h1e : _temp_cnt_T_159; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_161 = _temp_cnt_T_63[29] ? 6'h1d : _temp_cnt_T_160; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_162 = _temp_cnt_T_63[28] ? 6'h1c : _temp_cnt_T_161; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_163 = _temp_cnt_T_63[27] ? 6'h1b : _temp_cnt_T_162; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_164 = _temp_cnt_T_63[26] ? 6'h1a : _temp_cnt_T_163; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_165 = _temp_cnt_T_63[25] ? 6'h19 : _temp_cnt_T_164; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_166 = _temp_cnt_T_63[24] ? 6'h18 : _temp_cnt_T_165; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_167 = _temp_cnt_T_63[23] ? 6'h17 : _temp_cnt_T_166; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_168 = _temp_cnt_T_63[22] ? 6'h16 : _temp_cnt_T_167; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_169 = _temp_cnt_T_63[21] ? 6'h15 : _temp_cnt_T_168; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_170 = _temp_cnt_T_63[20] ? 6'h14 : _temp_cnt_T_169; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_171 = _temp_cnt_T_63[19] ? 6'h13 : _temp_cnt_T_170; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_172 = _temp_cnt_T_63[18] ? 6'h12 : _temp_cnt_T_171; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_173 = _temp_cnt_T_63[17] ? 6'h11 : _temp_cnt_T_172; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_174 = _temp_cnt_T_63[16] ? 6'h10 : _temp_cnt_T_173; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_175 = _temp_cnt_T_63[15] ? 6'hf : _temp_cnt_T_174; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_176 = _temp_cnt_T_63[14] ? 6'he : _temp_cnt_T_175; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_177 = _temp_cnt_T_63[13] ? 6'hd : _temp_cnt_T_176; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_178 = _temp_cnt_T_63[12] ? 6'hc : _temp_cnt_T_177; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_179 = _temp_cnt_T_63[11] ? 6'hb : _temp_cnt_T_178; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_180 = _temp_cnt_T_63[10] ? 6'ha : _temp_cnt_T_179; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_181 = _temp_cnt_T_63[9] ? 6'h9 : _temp_cnt_T_180; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_182 = _temp_cnt_T_63[8] ? 6'h8 : _temp_cnt_T_181; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_183 = _temp_cnt_T_63[7] ? 6'h7 : _temp_cnt_T_182; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_184 = _temp_cnt_T_63[6] ? 6'h6 : _temp_cnt_T_183; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_185 = _temp_cnt_T_63[5] ? 6'h5 : _temp_cnt_T_184; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_186 = _temp_cnt_T_63[4] ? 6'h4 : _temp_cnt_T_185; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_187 = _temp_cnt_T_63[3] ? 6'h3 : _temp_cnt_T_186; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_188 = _temp_cnt_T_63[2] ? 6'h2 : _temp_cnt_T_187; // @[Mux.scala 47:70]
  wire [5:0] _temp_cnt_T_189 = _temp_cnt_T_63[1] ? 6'h1 : _temp_cnt_T_188; // @[Mux.scala 47:70]
  wire [5:0] temp_cnt_1 = _temp_cnt_T_63[0] ? 6'h0 : _temp_cnt_T_189; // @[Mux.scala 47:70]
  wire [5:0] _io_cnt_T_1 = _temp_cnt_T_63[0] ? 6'h0 : _temp_cnt_T_189; // @[Cordic_LV.scala 110:32]
  wire [5:0] _io_cnt_T_4 = 6'sh0 - $signed(_io_cnt_T_1); // @[Cordic_LV.scala 110:15]
  wire [63:0] _io_out_T_1 = $signed(temp_x) >>> temp_cnt_1; // @[Cordic_LV.scala 111:23]
  wire [5:0] _GEN_98 = $signed(temp_x) > 64'sh100000000 ? $signed(_io_cnt_T_4) : $signed(6'sh0); // @[Cordic_LV.scala 110:12 113:12 98:78]
  wire [63:0] _GEN_99 = $signed(temp_x) > 64'sh100000000 ? $signed(_io_out_T_1) : $signed(temp_x); // @[Cordic_LV.scala 111:12 114:12 98:78]
  wire [94:0] _GEN_101 = $signed(temp_x) < 64'sh80000000 ? $signed(_io_out_T) : $signed({{31{_GEN_99[63]}},_GEN_99}); // @[Cordic_LV.scala 84:74 97:12]
  assign io_out = _GEN_101[63:0];
  assign io_cnt = $signed(temp_x) < 64'sh80000000 ? $signed({{1{_io_cnt_T[4]}},_io_cnt_T}) : $signed(_GEN_98); // @[Cordic_LV.scala 84:74 96:12]
  assign io_flag = $signed(io_x) < 64'sh0 ? 1'h0 : 1'h1; // @[Cordic_LV.scala 76:72 78:13 81:13]
endmodule
module CORDIC_LV_ORIGIN(
  input         clock,
  input         reset,
  input  [63:0] io_x,
  input  [63:0] io_y,
  output [63:0] io_z
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] current_x_0; // @[Cordic_LV.scala 25:43]
  reg [63:0] current_x_1; // @[Cordic_LV.scala 25:43]
  reg [63:0] current_x_2; // @[Cordic_LV.scala 25:43]
  reg [63:0] current_x_3; // @[Cordic_LV.scala 25:43]
  reg [63:0] current_x_4; // @[Cordic_LV.scala 25:43]
  reg [63:0] current_x_5; // @[Cordic_LV.scala 25:43]
  reg [63:0] current_x_6; // @[Cordic_LV.scala 25:43]
  reg [63:0] current_x_7; // @[Cordic_LV.scala 25:43]
  reg [63:0] current_x_8; // @[Cordic_LV.scala 25:43]
  reg [63:0] current_x_9; // @[Cordic_LV.scala 25:43]
  reg [63:0] current_x_10; // @[Cordic_LV.scala 25:43]
  reg [63:0] current_x_11; // @[Cordic_LV.scala 25:43]
  reg [63:0] current_x_12; // @[Cordic_LV.scala 25:43]
  reg [63:0] current_y_0; // @[Cordic_LV.scala 26:43]
  reg [63:0] current_y_1; // @[Cordic_LV.scala 26:43]
  reg [63:0] current_y_2; // @[Cordic_LV.scala 26:43]
  reg [63:0] current_y_3; // @[Cordic_LV.scala 26:43]
  reg [63:0] current_y_4; // @[Cordic_LV.scala 26:43]
  reg [63:0] current_y_5; // @[Cordic_LV.scala 26:43]
  reg [63:0] current_y_6; // @[Cordic_LV.scala 26:43]
  reg [63:0] current_y_7; // @[Cordic_LV.scala 26:43]
  reg [63:0] current_y_8; // @[Cordic_LV.scala 26:43]
  reg [63:0] current_y_9; // @[Cordic_LV.scala 26:43]
  reg [63:0] current_y_10; // @[Cordic_LV.scala 26:43]
  reg [63:0] current_y_11; // @[Cordic_LV.scala 26:43]
  reg [63:0] current_y_12; // @[Cordic_LV.scala 26:43]
  reg [63:0] current_y_13; // @[Cordic_LV.scala 26:43]
  reg [63:0] current_z_0; // @[Cordic_LV.scala 27:43]
  reg [63:0] current_z_1; // @[Cordic_LV.scala 27:43]
  reg [63:0] current_z_2; // @[Cordic_LV.scala 27:43]
  reg [63:0] current_z_3; // @[Cordic_LV.scala 27:43]
  reg [63:0] current_z_4; // @[Cordic_LV.scala 27:43]
  reg [63:0] current_z_5; // @[Cordic_LV.scala 27:43]
  reg [63:0] current_z_6; // @[Cordic_LV.scala 27:43]
  reg [63:0] current_z_7; // @[Cordic_LV.scala 27:43]
  reg [63:0] current_z_8; // @[Cordic_LV.scala 27:43]
  reg [63:0] current_z_9; // @[Cordic_LV.scala 27:43]
  reg [63:0] current_z_10; // @[Cordic_LV.scala 27:43]
  reg [63:0] current_z_11; // @[Cordic_LV.scala 27:43]
  reg [63:0] current_z_12; // @[Cordic_LV.scala 27:43]
  reg [63:0] current_z_13; // @[Cordic_LV.scala 27:43]
  reg [63:0] current_z_14; // @[Cordic_LV.scala 27:43]
  wire [63:0] _current_y_0_T_3 = $signed(io_y) - $signed(io_x); // @[Cordic_LV.scala 37:28]
  wire [62:0] _current_y_1_T = current_x_0[63:1]; // @[Cordic_LV.scala 42:62]
  wire [63:0] _GEN_28 = {{1{_current_y_1_T[62]}},_current_y_1_T}; // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_y_1_T_3 = $signed(current_y_0) + $signed(_GEN_28); // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_z_1_T_3 = $signed(current_z_0) - 64'sh80000000; // @[Cordic_LV.scala 43:42]
  wire [63:0] _current_y_1_T_7 = $signed(current_y_0) - $signed(_GEN_28); // @[Cordic_LV.scala 45:42]
  wire [63:0] _current_z_1_T_7 = $signed(current_z_0) + 64'sh80000000; // @[Cordic_LV.scala 46:42]
  wire [61:0] _current_y_2_T = current_x_1[63:2]; // @[Cordic_LV.scala 42:62]
  wire [63:0] _GEN_30 = {{2{_current_y_2_T[61]}},_current_y_2_T}; // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_y_2_T_3 = $signed(current_y_1) + $signed(_GEN_30); // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_z_2_T_3 = $signed(current_z_1) - 64'sh40000000; // @[Cordic_LV.scala 43:42]
  wire [63:0] _current_y_2_T_7 = $signed(current_y_1) - $signed(_GEN_30); // @[Cordic_LV.scala 45:42]
  wire [63:0] _current_z_2_T_7 = $signed(current_z_1) + 64'sh40000000; // @[Cordic_LV.scala 46:42]
  wire [60:0] _current_y_3_T = current_x_2[63:3]; // @[Cordic_LV.scala 42:62]
  wire [63:0] _GEN_32 = {{3{_current_y_3_T[60]}},_current_y_3_T}; // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_y_3_T_3 = $signed(current_y_2) + $signed(_GEN_32); // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_z_3_T_3 = $signed(current_z_2) - 64'sh20000000; // @[Cordic_LV.scala 43:42]
  wire [63:0] _current_y_3_T_7 = $signed(current_y_2) - $signed(_GEN_32); // @[Cordic_LV.scala 45:42]
  wire [63:0] _current_z_3_T_7 = $signed(current_z_2) + 64'sh20000000; // @[Cordic_LV.scala 46:42]
  wire [59:0] _current_y_4_T = current_x_3[63:4]; // @[Cordic_LV.scala 42:62]
  wire [63:0] _GEN_34 = {{4{_current_y_4_T[59]}},_current_y_4_T}; // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_y_4_T_3 = $signed(current_y_3) + $signed(_GEN_34); // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_z_4_T_3 = $signed(current_z_3) - 64'sh10000000; // @[Cordic_LV.scala 43:42]
  wire [63:0] _current_y_4_T_7 = $signed(current_y_3) - $signed(_GEN_34); // @[Cordic_LV.scala 45:42]
  wire [63:0] _current_z_4_T_7 = $signed(current_z_3) + 64'sh10000000; // @[Cordic_LV.scala 46:42]
  wire [58:0] _current_y_5_T = current_x_4[63:5]; // @[Cordic_LV.scala 42:62]
  wire [63:0] _GEN_36 = {{5{_current_y_5_T[58]}},_current_y_5_T}; // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_y_5_T_3 = $signed(current_y_4) + $signed(_GEN_36); // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_z_5_T_3 = $signed(current_z_4) - 64'sh8000000; // @[Cordic_LV.scala 43:42]
  wire [63:0] _current_y_5_T_7 = $signed(current_y_4) - $signed(_GEN_36); // @[Cordic_LV.scala 45:42]
  wire [63:0] _current_z_5_T_7 = $signed(current_z_4) + 64'sh8000000; // @[Cordic_LV.scala 46:42]
  wire [57:0] _current_y_6_T = current_x_5[63:6]; // @[Cordic_LV.scala 42:62]
  wire [63:0] _GEN_38 = {{6{_current_y_6_T[57]}},_current_y_6_T}; // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_y_6_T_3 = $signed(current_y_5) + $signed(_GEN_38); // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_z_6_T_3 = $signed(current_z_5) - 64'sh4000000; // @[Cordic_LV.scala 43:42]
  wire [63:0] _current_y_6_T_7 = $signed(current_y_5) - $signed(_GEN_38); // @[Cordic_LV.scala 45:42]
  wire [63:0] _current_z_6_T_7 = $signed(current_z_5) + 64'sh4000000; // @[Cordic_LV.scala 46:42]
  wire [56:0] _current_y_7_T = current_x_6[63:7]; // @[Cordic_LV.scala 42:62]
  wire [63:0] _GEN_40 = {{7{_current_y_7_T[56]}},_current_y_7_T}; // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_y_7_T_3 = $signed(current_y_6) + $signed(_GEN_40); // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_z_7_T_3 = $signed(current_z_6) - 64'sh2000000; // @[Cordic_LV.scala 43:42]
  wire [63:0] _current_y_7_T_7 = $signed(current_y_6) - $signed(_GEN_40); // @[Cordic_LV.scala 45:42]
  wire [63:0] _current_z_7_T_7 = $signed(current_z_6) + 64'sh2000000; // @[Cordic_LV.scala 46:42]
  wire [55:0] _current_y_8_T = current_x_7[63:8]; // @[Cordic_LV.scala 42:62]
  wire [63:0] _GEN_42 = {{8{_current_y_8_T[55]}},_current_y_8_T}; // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_y_8_T_3 = $signed(current_y_7) + $signed(_GEN_42); // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_z_8_T_3 = $signed(current_z_7) - 64'sh1000000; // @[Cordic_LV.scala 43:42]
  wire [63:0] _current_y_8_T_7 = $signed(current_y_7) - $signed(_GEN_42); // @[Cordic_LV.scala 45:42]
  wire [63:0] _current_z_8_T_7 = $signed(current_z_7) + 64'sh1000000; // @[Cordic_LV.scala 46:42]
  wire [54:0] _current_y_9_T = current_x_8[63:9]; // @[Cordic_LV.scala 42:62]
  wire [63:0] _GEN_44 = {{9{_current_y_9_T[54]}},_current_y_9_T}; // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_y_9_T_3 = $signed(current_y_8) + $signed(_GEN_44); // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_z_9_T_3 = $signed(current_z_8) - 64'sh800000; // @[Cordic_LV.scala 43:42]
  wire [63:0] _current_y_9_T_7 = $signed(current_y_8) - $signed(_GEN_44); // @[Cordic_LV.scala 45:42]
  wire [63:0] _current_z_9_T_7 = $signed(current_z_8) + 64'sh800000; // @[Cordic_LV.scala 46:42]
  wire [53:0] _current_y_10_T = current_x_9[63:10]; // @[Cordic_LV.scala 42:62]
  wire [63:0] _GEN_46 = {{10{_current_y_10_T[53]}},_current_y_10_T}; // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_y_10_T_3 = $signed(current_y_9) + $signed(_GEN_46); // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_z_10_T_3 = $signed(current_z_9) - 64'sh400000; // @[Cordic_LV.scala 43:42]
  wire [63:0] _current_y_10_T_7 = $signed(current_y_9) - $signed(_GEN_46); // @[Cordic_LV.scala 45:42]
  wire [63:0] _current_z_10_T_7 = $signed(current_z_9) + 64'sh400000; // @[Cordic_LV.scala 46:42]
  wire [52:0] _current_y_11_T = current_x_10[63:11]; // @[Cordic_LV.scala 42:62]
  wire [63:0] _GEN_48 = {{11{_current_y_11_T[52]}},_current_y_11_T}; // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_y_11_T_3 = $signed(current_y_10) + $signed(_GEN_48); // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_z_11_T_3 = $signed(current_z_10) - 64'sh200000; // @[Cordic_LV.scala 43:42]
  wire [63:0] _current_y_11_T_7 = $signed(current_y_10) - $signed(_GEN_48); // @[Cordic_LV.scala 45:42]
  wire [63:0] _current_z_11_T_7 = $signed(current_z_10) + 64'sh200000; // @[Cordic_LV.scala 46:42]
  wire [51:0] _current_y_12_T = current_x_11[63:12]; // @[Cordic_LV.scala 42:62]
  wire [63:0] _GEN_50 = {{12{_current_y_12_T[51]}},_current_y_12_T}; // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_y_12_T_3 = $signed(current_y_11) + $signed(_GEN_50); // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_z_12_T_3 = $signed(current_z_11) - 64'sh100000; // @[Cordic_LV.scala 43:42]
  wire [63:0] _current_y_12_T_7 = $signed(current_y_11) - $signed(_GEN_50); // @[Cordic_LV.scala 45:42]
  wire [63:0] _current_z_12_T_7 = $signed(current_z_11) + 64'sh100000; // @[Cordic_LV.scala 46:42]
  wire [50:0] _current_y_13_T = current_x_12[63:13]; // @[Cordic_LV.scala 42:62]
  wire [63:0] _GEN_52 = {{13{_current_y_13_T[50]}},_current_y_13_T}; // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_y_13_T_3 = $signed(current_y_12) + $signed(_GEN_52); // @[Cordic_LV.scala 42:42]
  wire [63:0] _current_z_13_T_3 = $signed(current_z_12) - 64'sh80000; // @[Cordic_LV.scala 43:42]
  wire [63:0] _current_y_13_T_7 = $signed(current_y_12) - $signed(_GEN_52); // @[Cordic_LV.scala 45:42]
  wire [63:0] _current_z_13_T_7 = $signed(current_z_12) + 64'sh80000; // @[Cordic_LV.scala 46:42]
  wire [63:0] _current_z_14_T_3 = $signed(current_z_13) - 64'sh40000; // @[Cordic_LV.scala 43:42]
  wire [63:0] _current_z_14_T_7 = $signed(current_z_13) + 64'sh40000; // @[Cordic_LV.scala 46:42]
  assign io_z = current_z_14; // @[Cordic_LV.scala 56:8]
  always @(posedge clock) begin
    if (reset) begin // @[Cordic_LV.scala 25:43]
      current_x_0 <= 64'sh0; // @[Cordic_LV.scala 25:43]
    end else begin
      current_x_0 <= io_x; // @[Cordic_LV.scala 36:20]
    end
    if (reset) begin // @[Cordic_LV.scala 25:43]
      current_x_1 <= 64'sh0; // @[Cordic_LV.scala 25:43]
    end else begin
      current_x_1 <= current_x_0; // @[Cordic_LV.scala 40:20]
    end
    if (reset) begin // @[Cordic_LV.scala 25:43]
      current_x_2 <= 64'sh0; // @[Cordic_LV.scala 25:43]
    end else begin
      current_x_2 <= current_x_1; // @[Cordic_LV.scala 40:20]
    end
    if (reset) begin // @[Cordic_LV.scala 25:43]
      current_x_3 <= 64'sh0; // @[Cordic_LV.scala 25:43]
    end else begin
      current_x_3 <= current_x_2; // @[Cordic_LV.scala 40:20]
    end
    if (reset) begin // @[Cordic_LV.scala 25:43]
      current_x_4 <= 64'sh0; // @[Cordic_LV.scala 25:43]
    end else begin
      current_x_4 <= current_x_3; // @[Cordic_LV.scala 40:20]
    end
    if (reset) begin // @[Cordic_LV.scala 25:43]
      current_x_5 <= 64'sh0; // @[Cordic_LV.scala 25:43]
    end else begin
      current_x_5 <= current_x_4; // @[Cordic_LV.scala 40:20]
    end
    if (reset) begin // @[Cordic_LV.scala 25:43]
      current_x_6 <= 64'sh0; // @[Cordic_LV.scala 25:43]
    end else begin
      current_x_6 <= current_x_5; // @[Cordic_LV.scala 40:20]
    end
    if (reset) begin // @[Cordic_LV.scala 25:43]
      current_x_7 <= 64'sh0; // @[Cordic_LV.scala 25:43]
    end else begin
      current_x_7 <= current_x_6; // @[Cordic_LV.scala 40:20]
    end
    if (reset) begin // @[Cordic_LV.scala 25:43]
      current_x_8 <= 64'sh0; // @[Cordic_LV.scala 25:43]
    end else begin
      current_x_8 <= current_x_7; // @[Cordic_LV.scala 40:20]
    end
    if (reset) begin // @[Cordic_LV.scala 25:43]
      current_x_9 <= 64'sh0; // @[Cordic_LV.scala 25:43]
    end else begin
      current_x_9 <= current_x_8; // @[Cordic_LV.scala 40:20]
    end
    if (reset) begin // @[Cordic_LV.scala 25:43]
      current_x_10 <= 64'sh0; // @[Cordic_LV.scala 25:43]
    end else begin
      current_x_10 <= current_x_9; // @[Cordic_LV.scala 40:20]
    end
    if (reset) begin // @[Cordic_LV.scala 25:43]
      current_x_11 <= 64'sh0; // @[Cordic_LV.scala 25:43]
    end else begin
      current_x_11 <= current_x_10; // @[Cordic_LV.scala 40:20]
    end
    if (reset) begin // @[Cordic_LV.scala 25:43]
      current_x_12 <= 64'sh0; // @[Cordic_LV.scala 25:43]
    end else begin
      current_x_12 <= current_x_11; // @[Cordic_LV.scala 40:20]
    end
    if (reset) begin // @[Cordic_LV.scala 26:43]
      current_y_0 <= 64'sh0; // @[Cordic_LV.scala 26:43]
    end else begin
      current_y_0 <= _current_y_0_T_3; // @[Cordic_LV.scala 37:20]
    end
    if (reset) begin // @[Cordic_LV.scala 26:43]
      current_y_1 <= 64'sh0; // @[Cordic_LV.scala 26:43]
    end else if ($signed(current_y_0) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_y_1 <= _current_y_1_T_3; // @[Cordic_LV.scala 42:22]
    end else begin
      current_y_1 <= _current_y_1_T_7; // @[Cordic_LV.scala 45:22]
    end
    if (reset) begin // @[Cordic_LV.scala 26:43]
      current_y_2 <= 64'sh0; // @[Cordic_LV.scala 26:43]
    end else if ($signed(current_y_1) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_y_2 <= _current_y_2_T_3; // @[Cordic_LV.scala 42:22]
    end else begin
      current_y_2 <= _current_y_2_T_7; // @[Cordic_LV.scala 45:22]
    end
    if (reset) begin // @[Cordic_LV.scala 26:43]
      current_y_3 <= 64'sh0; // @[Cordic_LV.scala 26:43]
    end else if ($signed(current_y_2) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_y_3 <= _current_y_3_T_3; // @[Cordic_LV.scala 42:22]
    end else begin
      current_y_3 <= _current_y_3_T_7; // @[Cordic_LV.scala 45:22]
    end
    if (reset) begin // @[Cordic_LV.scala 26:43]
      current_y_4 <= 64'sh0; // @[Cordic_LV.scala 26:43]
    end else if ($signed(current_y_3) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_y_4 <= _current_y_4_T_3; // @[Cordic_LV.scala 42:22]
    end else begin
      current_y_4 <= _current_y_4_T_7; // @[Cordic_LV.scala 45:22]
    end
    if (reset) begin // @[Cordic_LV.scala 26:43]
      current_y_5 <= 64'sh0; // @[Cordic_LV.scala 26:43]
    end else if ($signed(current_y_4) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_y_5 <= _current_y_5_T_3; // @[Cordic_LV.scala 42:22]
    end else begin
      current_y_5 <= _current_y_5_T_7; // @[Cordic_LV.scala 45:22]
    end
    if (reset) begin // @[Cordic_LV.scala 26:43]
      current_y_6 <= 64'sh0; // @[Cordic_LV.scala 26:43]
    end else if ($signed(current_y_5) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_y_6 <= _current_y_6_T_3; // @[Cordic_LV.scala 42:22]
    end else begin
      current_y_6 <= _current_y_6_T_7; // @[Cordic_LV.scala 45:22]
    end
    if (reset) begin // @[Cordic_LV.scala 26:43]
      current_y_7 <= 64'sh0; // @[Cordic_LV.scala 26:43]
    end else if ($signed(current_y_6) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_y_7 <= _current_y_7_T_3; // @[Cordic_LV.scala 42:22]
    end else begin
      current_y_7 <= _current_y_7_T_7; // @[Cordic_LV.scala 45:22]
    end
    if (reset) begin // @[Cordic_LV.scala 26:43]
      current_y_8 <= 64'sh0; // @[Cordic_LV.scala 26:43]
    end else if ($signed(current_y_7) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_y_8 <= _current_y_8_T_3; // @[Cordic_LV.scala 42:22]
    end else begin
      current_y_8 <= _current_y_8_T_7; // @[Cordic_LV.scala 45:22]
    end
    if (reset) begin // @[Cordic_LV.scala 26:43]
      current_y_9 <= 64'sh0; // @[Cordic_LV.scala 26:43]
    end else if ($signed(current_y_8) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_y_9 <= _current_y_9_T_3; // @[Cordic_LV.scala 42:22]
    end else begin
      current_y_9 <= _current_y_9_T_7; // @[Cordic_LV.scala 45:22]
    end
    if (reset) begin // @[Cordic_LV.scala 26:43]
      current_y_10 <= 64'sh0; // @[Cordic_LV.scala 26:43]
    end else if ($signed(current_y_9) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_y_10 <= _current_y_10_T_3; // @[Cordic_LV.scala 42:22]
    end else begin
      current_y_10 <= _current_y_10_T_7; // @[Cordic_LV.scala 45:22]
    end
    if (reset) begin // @[Cordic_LV.scala 26:43]
      current_y_11 <= 64'sh0; // @[Cordic_LV.scala 26:43]
    end else if ($signed(current_y_10) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_y_11 <= _current_y_11_T_3; // @[Cordic_LV.scala 42:22]
    end else begin
      current_y_11 <= _current_y_11_T_7; // @[Cordic_LV.scala 45:22]
    end
    if (reset) begin // @[Cordic_LV.scala 26:43]
      current_y_12 <= 64'sh0; // @[Cordic_LV.scala 26:43]
    end else if ($signed(current_y_11) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_y_12 <= _current_y_12_T_3; // @[Cordic_LV.scala 42:22]
    end else begin
      current_y_12 <= _current_y_12_T_7; // @[Cordic_LV.scala 45:22]
    end
    if (reset) begin // @[Cordic_LV.scala 26:43]
      current_y_13 <= 64'sh0; // @[Cordic_LV.scala 26:43]
    end else if ($signed(current_y_12) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_y_13 <= _current_y_13_T_3; // @[Cordic_LV.scala 42:22]
    end else begin
      current_y_13 <= _current_y_13_T_7; // @[Cordic_LV.scala 45:22]
    end
    if (reset) begin // @[Cordic_LV.scala 27:43]
      current_z_0 <= 64'sh0; // @[Cordic_LV.scala 27:43]
    end else begin
      current_z_0 <= 64'sh100000000; // @[Cordic_LV.scala 38:20]
    end
    if (reset) begin // @[Cordic_LV.scala 27:43]
      current_z_1 <= 64'sh0; // @[Cordic_LV.scala 27:43]
    end else if ($signed(current_y_0) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_z_1 <= _current_z_1_T_3; // @[Cordic_LV.scala 43:22]
    end else begin
      current_z_1 <= _current_z_1_T_7; // @[Cordic_LV.scala 46:22]
    end
    if (reset) begin // @[Cordic_LV.scala 27:43]
      current_z_2 <= 64'sh0; // @[Cordic_LV.scala 27:43]
    end else if ($signed(current_y_1) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_z_2 <= _current_z_2_T_3; // @[Cordic_LV.scala 43:22]
    end else begin
      current_z_2 <= _current_z_2_T_7; // @[Cordic_LV.scala 46:22]
    end
    if (reset) begin // @[Cordic_LV.scala 27:43]
      current_z_3 <= 64'sh0; // @[Cordic_LV.scala 27:43]
    end else if ($signed(current_y_2) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_z_3 <= _current_z_3_T_3; // @[Cordic_LV.scala 43:22]
    end else begin
      current_z_3 <= _current_z_3_T_7; // @[Cordic_LV.scala 46:22]
    end
    if (reset) begin // @[Cordic_LV.scala 27:43]
      current_z_4 <= 64'sh0; // @[Cordic_LV.scala 27:43]
    end else if ($signed(current_y_3) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_z_4 <= _current_z_4_T_3; // @[Cordic_LV.scala 43:22]
    end else begin
      current_z_4 <= _current_z_4_T_7; // @[Cordic_LV.scala 46:22]
    end
    if (reset) begin // @[Cordic_LV.scala 27:43]
      current_z_5 <= 64'sh0; // @[Cordic_LV.scala 27:43]
    end else if ($signed(current_y_4) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_z_5 <= _current_z_5_T_3; // @[Cordic_LV.scala 43:22]
    end else begin
      current_z_5 <= _current_z_5_T_7; // @[Cordic_LV.scala 46:22]
    end
    if (reset) begin // @[Cordic_LV.scala 27:43]
      current_z_6 <= 64'sh0; // @[Cordic_LV.scala 27:43]
    end else if ($signed(current_y_5) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_z_6 <= _current_z_6_T_3; // @[Cordic_LV.scala 43:22]
    end else begin
      current_z_6 <= _current_z_6_T_7; // @[Cordic_LV.scala 46:22]
    end
    if (reset) begin // @[Cordic_LV.scala 27:43]
      current_z_7 <= 64'sh0; // @[Cordic_LV.scala 27:43]
    end else if ($signed(current_y_6) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_z_7 <= _current_z_7_T_3; // @[Cordic_LV.scala 43:22]
    end else begin
      current_z_7 <= _current_z_7_T_7; // @[Cordic_LV.scala 46:22]
    end
    if (reset) begin // @[Cordic_LV.scala 27:43]
      current_z_8 <= 64'sh0; // @[Cordic_LV.scala 27:43]
    end else if ($signed(current_y_7) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_z_8 <= _current_z_8_T_3; // @[Cordic_LV.scala 43:22]
    end else begin
      current_z_8 <= _current_z_8_T_7; // @[Cordic_LV.scala 46:22]
    end
    if (reset) begin // @[Cordic_LV.scala 27:43]
      current_z_9 <= 64'sh0; // @[Cordic_LV.scala 27:43]
    end else if ($signed(current_y_8) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_z_9 <= _current_z_9_T_3; // @[Cordic_LV.scala 43:22]
    end else begin
      current_z_9 <= _current_z_9_T_7; // @[Cordic_LV.scala 46:22]
    end
    if (reset) begin // @[Cordic_LV.scala 27:43]
      current_z_10 <= 64'sh0; // @[Cordic_LV.scala 27:43]
    end else if ($signed(current_y_9) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_z_10 <= _current_z_10_T_3; // @[Cordic_LV.scala 43:22]
    end else begin
      current_z_10 <= _current_z_10_T_7; // @[Cordic_LV.scala 46:22]
    end
    if (reset) begin // @[Cordic_LV.scala 27:43]
      current_z_11 <= 64'sh0; // @[Cordic_LV.scala 27:43]
    end else if ($signed(current_y_10) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_z_11 <= _current_z_11_T_3; // @[Cordic_LV.scala 43:22]
    end else begin
      current_z_11 <= _current_z_11_T_7; // @[Cordic_LV.scala 46:22]
    end
    if (reset) begin // @[Cordic_LV.scala 27:43]
      current_z_12 <= 64'sh0; // @[Cordic_LV.scala 27:43]
    end else if ($signed(current_y_11) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_z_12 <= _current_z_12_T_3; // @[Cordic_LV.scala 43:22]
    end else begin
      current_z_12 <= _current_z_12_T_7; // @[Cordic_LV.scala 46:22]
    end
    if (reset) begin // @[Cordic_LV.scala 27:43]
      current_z_13 <= 64'sh0; // @[Cordic_LV.scala 27:43]
    end else if ($signed(current_y_12) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_z_13 <= _current_z_13_T_3; // @[Cordic_LV.scala 43:22]
    end else begin
      current_z_13 <= _current_z_13_T_7; // @[Cordic_LV.scala 46:22]
    end
    if (reset) begin // @[Cordic_LV.scala 27:43]
      current_z_14 <= 64'sh0; // @[Cordic_LV.scala 27:43]
    end else if ($signed(current_y_13) < 64'sh0) begin // @[Cordic_LV.scala 41:88]
      current_z_14 <= _current_z_14_T_3; // @[Cordic_LV.scala 43:22]
    end else begin
      current_z_14 <= _current_z_14_T_7; // @[Cordic_LV.scala 46:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  current_x_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  current_x_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  current_x_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  current_x_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  current_x_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  current_x_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  current_x_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  current_x_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  current_x_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  current_x_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  current_x_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  current_x_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  current_x_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  current_y_0 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  current_y_1 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  current_y_2 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  current_y_3 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  current_y_4 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  current_y_5 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  current_y_6 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  current_y_7 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  current_y_8 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  current_y_9 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  current_y_10 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  current_y_11 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  current_y_12 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  current_y_13 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  current_z_0 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  current_z_1 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  current_z_2 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  current_z_3 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  current_z_4 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  current_z_5 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  current_z_6 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  current_z_7 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  current_z_8 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  current_z_9 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  current_z_10 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  current_z_11 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  current_z_12 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  current_z_13 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  current_z_14 = _RAND_41[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cordic_divide(
  input         clock,
  input         reset,
  input  [63:0] io_x,
  input  [63:0] io_y,
  output [63:0] io_z
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] unit_io_x; // @[Cordic_LV.scala 131:22]
  wire [63:0] unit_io_out; // @[Cordic_LV.scala 131:22]
  wire [5:0] unit_io_cnt; // @[Cordic_LV.scala 131:22]
  wire  unit_io_flag; // @[Cordic_LV.scala 131:22]
  wire [63:0] unit_1_io_x; // @[Cordic_LV.scala 131:22]
  wire [63:0] unit_1_io_out; // @[Cordic_LV.scala 131:22]
  wire [5:0] unit_1_io_cnt; // @[Cordic_LV.scala 131:22]
  wire  unit_1_io_flag; // @[Cordic_LV.scala 131:22]
  wire  cordic_lv_clock; // @[Cordic_LV.scala 177:43]
  wire  cordic_lv_reset; // @[Cordic_LV.scala 177:43]
  wire [63:0] cordic_lv_io_x; // @[Cordic_LV.scala 177:43]
  wire [63:0] cordic_lv_io_y; // @[Cordic_LV.scala 177:43]
  wire [63:0] cordic_lv_io_z; // @[Cordic_LV.scala 177:43]
  reg [5:0] x_cnt_reg_0; // @[Cordic_LV.scala 158:37]
  reg [5:0] x_cnt_reg_1; // @[Cordic_LV.scala 158:37]
  reg [5:0] x_cnt_reg_2; // @[Cordic_LV.scala 158:37]
  reg [5:0] x_cnt_reg_3; // @[Cordic_LV.scala 158:37]
  reg [5:0] x_cnt_reg_4; // @[Cordic_LV.scala 158:37]
  reg [5:0] x_cnt_reg_5; // @[Cordic_LV.scala 158:37]
  reg [5:0] x_cnt_reg_6; // @[Cordic_LV.scala 158:37]
  reg [5:0] x_cnt_reg_7; // @[Cordic_LV.scala 158:37]
  reg [5:0] x_cnt_reg_8; // @[Cordic_LV.scala 158:37]
  reg [5:0] x_cnt_reg_9; // @[Cordic_LV.scala 158:37]
  reg [5:0] x_cnt_reg_10; // @[Cordic_LV.scala 158:37]
  reg [5:0] x_cnt_reg_11; // @[Cordic_LV.scala 158:37]
  reg [5:0] x_cnt_reg_12; // @[Cordic_LV.scala 158:37]
  reg [5:0] x_cnt_reg_13; // @[Cordic_LV.scala 158:37]
  reg [5:0] x_cnt_reg_14; // @[Cordic_LV.scala 158:37]
  reg  x_flag_reg_0; // @[Cordic_LV.scala 159:38]
  reg  x_flag_reg_1; // @[Cordic_LV.scala 159:38]
  reg  x_flag_reg_2; // @[Cordic_LV.scala 159:38]
  reg  x_flag_reg_3; // @[Cordic_LV.scala 159:38]
  reg  x_flag_reg_4; // @[Cordic_LV.scala 159:38]
  reg  x_flag_reg_5; // @[Cordic_LV.scala 159:38]
  reg  x_flag_reg_6; // @[Cordic_LV.scala 159:38]
  reg  x_flag_reg_7; // @[Cordic_LV.scala 159:38]
  reg  x_flag_reg_8; // @[Cordic_LV.scala 159:38]
  reg  x_flag_reg_9; // @[Cordic_LV.scala 159:38]
  reg  x_flag_reg_10; // @[Cordic_LV.scala 159:38]
  reg  x_flag_reg_11; // @[Cordic_LV.scala 159:38]
  reg  x_flag_reg_12; // @[Cordic_LV.scala 159:38]
  reg  x_flag_reg_13; // @[Cordic_LV.scala 159:38]
  reg  x_flag_reg_14; // @[Cordic_LV.scala 159:38]
  reg [5:0] y_cnt_reg_0; // @[Cordic_LV.scala 160:37]
  reg [5:0] y_cnt_reg_1; // @[Cordic_LV.scala 160:37]
  reg [5:0] y_cnt_reg_2; // @[Cordic_LV.scala 160:37]
  reg [5:0] y_cnt_reg_3; // @[Cordic_LV.scala 160:37]
  reg [5:0] y_cnt_reg_4; // @[Cordic_LV.scala 160:37]
  reg [5:0] y_cnt_reg_5; // @[Cordic_LV.scala 160:37]
  reg [5:0] y_cnt_reg_6; // @[Cordic_LV.scala 160:37]
  reg [5:0] y_cnt_reg_7; // @[Cordic_LV.scala 160:37]
  reg [5:0] y_cnt_reg_8; // @[Cordic_LV.scala 160:37]
  reg [5:0] y_cnt_reg_9; // @[Cordic_LV.scala 160:37]
  reg [5:0] y_cnt_reg_10; // @[Cordic_LV.scala 160:37]
  reg [5:0] y_cnt_reg_11; // @[Cordic_LV.scala 160:37]
  reg [5:0] y_cnt_reg_12; // @[Cordic_LV.scala 160:37]
  reg [5:0] y_cnt_reg_13; // @[Cordic_LV.scala 160:37]
  reg [5:0] y_cnt_reg_14; // @[Cordic_LV.scala 160:37]
  reg  y_flag_reg_0; // @[Cordic_LV.scala 161:38]
  reg  y_flag_reg_1; // @[Cordic_LV.scala 161:38]
  reg  y_flag_reg_2; // @[Cordic_LV.scala 161:38]
  reg  y_flag_reg_3; // @[Cordic_LV.scala 161:38]
  reg  y_flag_reg_4; // @[Cordic_LV.scala 161:38]
  reg  y_flag_reg_5; // @[Cordic_LV.scala 161:38]
  reg  y_flag_reg_6; // @[Cordic_LV.scala 161:38]
  reg  y_flag_reg_7; // @[Cordic_LV.scala 161:38]
  reg  y_flag_reg_8; // @[Cordic_LV.scala 161:38]
  reg  y_flag_reg_9; // @[Cordic_LV.scala 161:38]
  reg  y_flag_reg_10; // @[Cordic_LV.scala 161:38]
  reg  y_flag_reg_11; // @[Cordic_LV.scala 161:38]
  reg  y_flag_reg_12; // @[Cordic_LV.scala 161:38]
  reg  y_flag_reg_13; // @[Cordic_LV.scala 161:38]
  reg  y_flag_reg_14; // @[Cordic_LV.scala 161:38]
  wire  _T_2 = x_flag_reg_14 & ~y_flag_reg_14; // @[Cordic_LV.scala 183:50]
  wire [63:0] _unnormed_z_T_2 = 64'sh0 - $signed(cordic_lv_io_z); // @[Cordic_LV.scala 185:19]
  wire [63:0] unnormed_z = _T_2 | ~x_flag_reg_14 & y_flag_reg_14 ? $signed(_unnormed_z_T_2) : $signed(cordic_lv_io_z); // @[Cordic_LV.scala 184:96 185:16 187:16]
  wire [5:0] shift_cnt = $signed(y_cnt_reg_14) - $signed(x_cnt_reg_14); // @[Cordic_LV.scala 189:49]
  wire [5:0] _io_z_T_3 = 6'sh0 - $signed(shift_cnt); // @[Cordic_LV.scala 191:46]
  wire [126:0] _GEN_0 = {{63{unnormed_z[63]}},unnormed_z}; // @[Cordic_LV.scala 191:24]
  wire [126:0] _io_z_T_4 = $signed(_GEN_0) << _io_z_T_3; // @[Cordic_LV.scala 191:24]
  wire [5:0] _io_z_T_5 = $signed(y_cnt_reg_14) - $signed(x_cnt_reg_14); // @[Cordic_LV.scala 193:43]
  wire [63:0] _io_z_T_6 = $signed(unnormed_z) >>> _io_z_T_5; // @[Cordic_LV.scala 193:24]
  wire [126:0] _GEN_1 = $signed(shift_cnt) < 6'sh0 ? $signed(_io_z_T_4) : $signed({{63{_io_z_T_6[63]}},_io_z_T_6}); // @[Cordic_LV.scala 190:25 191:10 193:10]
  shift_2_range unit ( // @[Cordic_LV.scala 131:22]
    .io_x(unit_io_x),
    .io_out(unit_io_out),
    .io_cnt(unit_io_cnt),
    .io_flag(unit_io_flag)
  );
  shift_2_range unit_1 ( // @[Cordic_LV.scala 131:22]
    .io_x(unit_1_io_x),
    .io_out(unit_1_io_out),
    .io_cnt(unit_1_io_cnt),
    .io_flag(unit_1_io_flag)
  );
  CORDIC_LV_ORIGIN cordic_lv ( // @[Cordic_LV.scala 177:43]
    .clock(cordic_lv_clock),
    .reset(cordic_lv_reset),
    .io_x(cordic_lv_io_x),
    .io_y(cordic_lv_io_y),
    .io_z(cordic_lv_io_z)
  );
  assign io_z = _GEN_1[63:0];
  assign unit_io_x = io_x; // @[Cordic_LV.scala 132:15]
  assign unit_1_io_x = io_y; // @[Cordic_LV.scala 132:15]
  assign cordic_lv_clock = clock;
  assign cordic_lv_reset = reset;
  assign cordic_lv_io_x = unit_io_out; // @[Cordic_LV.scala 178:18]
  assign cordic_lv_io_y = unit_1_io_out; // @[Cordic_LV.scala 179:18]
  always @(posedge clock) begin
    if (reset) begin // @[Cordic_LV.scala 158:37]
      x_cnt_reg_0 <= 6'sh0; // @[Cordic_LV.scala 158:37]
    end else begin
      x_cnt_reg_0 <= unit_io_cnt; // @[Cordic_LV.scala 164:20]
    end
    if (reset) begin // @[Cordic_LV.scala 158:37]
      x_cnt_reg_1 <= 6'sh0; // @[Cordic_LV.scala 158:37]
    end else begin
      x_cnt_reg_1 <= x_cnt_reg_0; // @[Cordic_LV.scala 169:20]
    end
    if (reset) begin // @[Cordic_LV.scala 158:37]
      x_cnt_reg_2 <= 6'sh0; // @[Cordic_LV.scala 158:37]
    end else begin
      x_cnt_reg_2 <= x_cnt_reg_1; // @[Cordic_LV.scala 169:20]
    end
    if (reset) begin // @[Cordic_LV.scala 158:37]
      x_cnt_reg_3 <= 6'sh0; // @[Cordic_LV.scala 158:37]
    end else begin
      x_cnt_reg_3 <= x_cnt_reg_2; // @[Cordic_LV.scala 169:20]
    end
    if (reset) begin // @[Cordic_LV.scala 158:37]
      x_cnt_reg_4 <= 6'sh0; // @[Cordic_LV.scala 158:37]
    end else begin
      x_cnt_reg_4 <= x_cnt_reg_3; // @[Cordic_LV.scala 169:20]
    end
    if (reset) begin // @[Cordic_LV.scala 158:37]
      x_cnt_reg_5 <= 6'sh0; // @[Cordic_LV.scala 158:37]
    end else begin
      x_cnt_reg_5 <= x_cnt_reg_4; // @[Cordic_LV.scala 169:20]
    end
    if (reset) begin // @[Cordic_LV.scala 158:37]
      x_cnt_reg_6 <= 6'sh0; // @[Cordic_LV.scala 158:37]
    end else begin
      x_cnt_reg_6 <= x_cnt_reg_5; // @[Cordic_LV.scala 169:20]
    end
    if (reset) begin // @[Cordic_LV.scala 158:37]
      x_cnt_reg_7 <= 6'sh0; // @[Cordic_LV.scala 158:37]
    end else begin
      x_cnt_reg_7 <= x_cnt_reg_6; // @[Cordic_LV.scala 169:20]
    end
    if (reset) begin // @[Cordic_LV.scala 158:37]
      x_cnt_reg_8 <= 6'sh0; // @[Cordic_LV.scala 158:37]
    end else begin
      x_cnt_reg_8 <= x_cnt_reg_7; // @[Cordic_LV.scala 169:20]
    end
    if (reset) begin // @[Cordic_LV.scala 158:37]
      x_cnt_reg_9 <= 6'sh0; // @[Cordic_LV.scala 158:37]
    end else begin
      x_cnt_reg_9 <= x_cnt_reg_8; // @[Cordic_LV.scala 169:20]
    end
    if (reset) begin // @[Cordic_LV.scala 158:37]
      x_cnt_reg_10 <= 6'sh0; // @[Cordic_LV.scala 158:37]
    end else begin
      x_cnt_reg_10 <= x_cnt_reg_9; // @[Cordic_LV.scala 169:20]
    end
    if (reset) begin // @[Cordic_LV.scala 158:37]
      x_cnt_reg_11 <= 6'sh0; // @[Cordic_LV.scala 158:37]
    end else begin
      x_cnt_reg_11 <= x_cnt_reg_10; // @[Cordic_LV.scala 169:20]
    end
    if (reset) begin // @[Cordic_LV.scala 158:37]
      x_cnt_reg_12 <= 6'sh0; // @[Cordic_LV.scala 158:37]
    end else begin
      x_cnt_reg_12 <= x_cnt_reg_11; // @[Cordic_LV.scala 169:20]
    end
    if (reset) begin // @[Cordic_LV.scala 158:37]
      x_cnt_reg_13 <= 6'sh0; // @[Cordic_LV.scala 158:37]
    end else begin
      x_cnt_reg_13 <= x_cnt_reg_12; // @[Cordic_LV.scala 169:20]
    end
    if (reset) begin // @[Cordic_LV.scala 158:37]
      x_cnt_reg_14 <= 6'sh0; // @[Cordic_LV.scala 158:37]
    end else begin
      x_cnt_reg_14 <= x_cnt_reg_13; // @[Cordic_LV.scala 169:20]
    end
    if (reset) begin // @[Cordic_LV.scala 159:38]
      x_flag_reg_0 <= 1'h0; // @[Cordic_LV.scala 159:38]
    end else begin
      x_flag_reg_0 <= unit_io_flag; // @[Cordic_LV.scala 165:21]
    end
    if (reset) begin // @[Cordic_LV.scala 159:38]
      x_flag_reg_1 <= 1'h0; // @[Cordic_LV.scala 159:38]
    end else begin
      x_flag_reg_1 <= x_flag_reg_0; // @[Cordic_LV.scala 170:21]
    end
    if (reset) begin // @[Cordic_LV.scala 159:38]
      x_flag_reg_2 <= 1'h0; // @[Cordic_LV.scala 159:38]
    end else begin
      x_flag_reg_2 <= x_flag_reg_1; // @[Cordic_LV.scala 170:21]
    end
    if (reset) begin // @[Cordic_LV.scala 159:38]
      x_flag_reg_3 <= 1'h0; // @[Cordic_LV.scala 159:38]
    end else begin
      x_flag_reg_3 <= x_flag_reg_2; // @[Cordic_LV.scala 170:21]
    end
    if (reset) begin // @[Cordic_LV.scala 159:38]
      x_flag_reg_4 <= 1'h0; // @[Cordic_LV.scala 159:38]
    end else begin
      x_flag_reg_4 <= x_flag_reg_3; // @[Cordic_LV.scala 170:21]
    end
    if (reset) begin // @[Cordic_LV.scala 159:38]
      x_flag_reg_5 <= 1'h0; // @[Cordic_LV.scala 159:38]
    end else begin
      x_flag_reg_5 <= x_flag_reg_4; // @[Cordic_LV.scala 170:21]
    end
    if (reset) begin // @[Cordic_LV.scala 159:38]
      x_flag_reg_6 <= 1'h0; // @[Cordic_LV.scala 159:38]
    end else begin
      x_flag_reg_6 <= x_flag_reg_5; // @[Cordic_LV.scala 170:21]
    end
    if (reset) begin // @[Cordic_LV.scala 159:38]
      x_flag_reg_7 <= 1'h0; // @[Cordic_LV.scala 159:38]
    end else begin
      x_flag_reg_7 <= x_flag_reg_6; // @[Cordic_LV.scala 170:21]
    end
    if (reset) begin // @[Cordic_LV.scala 159:38]
      x_flag_reg_8 <= 1'h0; // @[Cordic_LV.scala 159:38]
    end else begin
      x_flag_reg_8 <= x_flag_reg_7; // @[Cordic_LV.scala 170:21]
    end
    if (reset) begin // @[Cordic_LV.scala 159:38]
      x_flag_reg_9 <= 1'h0; // @[Cordic_LV.scala 159:38]
    end else begin
      x_flag_reg_9 <= x_flag_reg_8; // @[Cordic_LV.scala 170:21]
    end
    if (reset) begin // @[Cordic_LV.scala 159:38]
      x_flag_reg_10 <= 1'h0; // @[Cordic_LV.scala 159:38]
    end else begin
      x_flag_reg_10 <= x_flag_reg_9; // @[Cordic_LV.scala 170:21]
    end
    if (reset) begin // @[Cordic_LV.scala 159:38]
      x_flag_reg_11 <= 1'h0; // @[Cordic_LV.scala 159:38]
    end else begin
      x_flag_reg_11 <= x_flag_reg_10; // @[Cordic_LV.scala 170:21]
    end
    if (reset) begin // @[Cordic_LV.scala 159:38]
      x_flag_reg_12 <= 1'h0; // @[Cordic_LV.scala 159:38]
    end else begin
      x_flag_reg_12 <= x_flag_reg_11; // @[Cordic_LV.scala 170:21]
    end
    if (reset) begin // @[Cordic_LV.scala 159:38]
      x_flag_reg_13 <= 1'h0; // @[Cordic_LV.scala 159:38]
    end else begin
      x_flag_reg_13 <= x_flag_reg_12; // @[Cordic_LV.scala 170:21]
    end
    if (reset) begin // @[Cordic_LV.scala 159:38]
      x_flag_reg_14 <= 1'h0; // @[Cordic_LV.scala 159:38]
    end else begin
      x_flag_reg_14 <= x_flag_reg_13; // @[Cordic_LV.scala 170:21]
    end
    if (reset) begin // @[Cordic_LV.scala 160:37]
      y_cnt_reg_0 <= 6'sh0; // @[Cordic_LV.scala 160:37]
    end else begin
      y_cnt_reg_0 <= unit_1_io_cnt; // @[Cordic_LV.scala 166:20]
    end
    if (reset) begin // @[Cordic_LV.scala 160:37]
      y_cnt_reg_1 <= 6'sh0; // @[Cordic_LV.scala 160:37]
    end else begin
      y_cnt_reg_1 <= y_cnt_reg_0; // @[Cordic_LV.scala 171:20]
    end
    if (reset) begin // @[Cordic_LV.scala 160:37]
      y_cnt_reg_2 <= 6'sh0; // @[Cordic_LV.scala 160:37]
    end else begin
      y_cnt_reg_2 <= y_cnt_reg_1; // @[Cordic_LV.scala 171:20]
    end
    if (reset) begin // @[Cordic_LV.scala 160:37]
      y_cnt_reg_3 <= 6'sh0; // @[Cordic_LV.scala 160:37]
    end else begin
      y_cnt_reg_3 <= y_cnt_reg_2; // @[Cordic_LV.scala 171:20]
    end
    if (reset) begin // @[Cordic_LV.scala 160:37]
      y_cnt_reg_4 <= 6'sh0; // @[Cordic_LV.scala 160:37]
    end else begin
      y_cnt_reg_4 <= y_cnt_reg_3; // @[Cordic_LV.scala 171:20]
    end
    if (reset) begin // @[Cordic_LV.scala 160:37]
      y_cnt_reg_5 <= 6'sh0; // @[Cordic_LV.scala 160:37]
    end else begin
      y_cnt_reg_5 <= y_cnt_reg_4; // @[Cordic_LV.scala 171:20]
    end
    if (reset) begin // @[Cordic_LV.scala 160:37]
      y_cnt_reg_6 <= 6'sh0; // @[Cordic_LV.scala 160:37]
    end else begin
      y_cnt_reg_6 <= y_cnt_reg_5; // @[Cordic_LV.scala 171:20]
    end
    if (reset) begin // @[Cordic_LV.scala 160:37]
      y_cnt_reg_7 <= 6'sh0; // @[Cordic_LV.scala 160:37]
    end else begin
      y_cnt_reg_7 <= y_cnt_reg_6; // @[Cordic_LV.scala 171:20]
    end
    if (reset) begin // @[Cordic_LV.scala 160:37]
      y_cnt_reg_8 <= 6'sh0; // @[Cordic_LV.scala 160:37]
    end else begin
      y_cnt_reg_8 <= y_cnt_reg_7; // @[Cordic_LV.scala 171:20]
    end
    if (reset) begin // @[Cordic_LV.scala 160:37]
      y_cnt_reg_9 <= 6'sh0; // @[Cordic_LV.scala 160:37]
    end else begin
      y_cnt_reg_9 <= y_cnt_reg_8; // @[Cordic_LV.scala 171:20]
    end
    if (reset) begin // @[Cordic_LV.scala 160:37]
      y_cnt_reg_10 <= 6'sh0; // @[Cordic_LV.scala 160:37]
    end else begin
      y_cnt_reg_10 <= y_cnt_reg_9; // @[Cordic_LV.scala 171:20]
    end
    if (reset) begin // @[Cordic_LV.scala 160:37]
      y_cnt_reg_11 <= 6'sh0; // @[Cordic_LV.scala 160:37]
    end else begin
      y_cnt_reg_11 <= y_cnt_reg_10; // @[Cordic_LV.scala 171:20]
    end
    if (reset) begin // @[Cordic_LV.scala 160:37]
      y_cnt_reg_12 <= 6'sh0; // @[Cordic_LV.scala 160:37]
    end else begin
      y_cnt_reg_12 <= y_cnt_reg_11; // @[Cordic_LV.scala 171:20]
    end
    if (reset) begin // @[Cordic_LV.scala 160:37]
      y_cnt_reg_13 <= 6'sh0; // @[Cordic_LV.scala 160:37]
    end else begin
      y_cnt_reg_13 <= y_cnt_reg_12; // @[Cordic_LV.scala 171:20]
    end
    if (reset) begin // @[Cordic_LV.scala 160:37]
      y_cnt_reg_14 <= 6'sh0; // @[Cordic_LV.scala 160:37]
    end else begin
      y_cnt_reg_14 <= y_cnt_reg_13; // @[Cordic_LV.scala 171:20]
    end
    if (reset) begin // @[Cordic_LV.scala 161:38]
      y_flag_reg_0 <= 1'h0; // @[Cordic_LV.scala 161:38]
    end else begin
      y_flag_reg_0 <= unit_1_io_flag; // @[Cordic_LV.scala 167:21]
    end
    if (reset) begin // @[Cordic_LV.scala 161:38]
      y_flag_reg_1 <= 1'h0; // @[Cordic_LV.scala 161:38]
    end else begin
      y_flag_reg_1 <= y_flag_reg_0; // @[Cordic_LV.scala 172:21]
    end
    if (reset) begin // @[Cordic_LV.scala 161:38]
      y_flag_reg_2 <= 1'h0; // @[Cordic_LV.scala 161:38]
    end else begin
      y_flag_reg_2 <= y_flag_reg_1; // @[Cordic_LV.scala 172:21]
    end
    if (reset) begin // @[Cordic_LV.scala 161:38]
      y_flag_reg_3 <= 1'h0; // @[Cordic_LV.scala 161:38]
    end else begin
      y_flag_reg_3 <= y_flag_reg_2; // @[Cordic_LV.scala 172:21]
    end
    if (reset) begin // @[Cordic_LV.scala 161:38]
      y_flag_reg_4 <= 1'h0; // @[Cordic_LV.scala 161:38]
    end else begin
      y_flag_reg_4 <= y_flag_reg_3; // @[Cordic_LV.scala 172:21]
    end
    if (reset) begin // @[Cordic_LV.scala 161:38]
      y_flag_reg_5 <= 1'h0; // @[Cordic_LV.scala 161:38]
    end else begin
      y_flag_reg_5 <= y_flag_reg_4; // @[Cordic_LV.scala 172:21]
    end
    if (reset) begin // @[Cordic_LV.scala 161:38]
      y_flag_reg_6 <= 1'h0; // @[Cordic_LV.scala 161:38]
    end else begin
      y_flag_reg_6 <= y_flag_reg_5; // @[Cordic_LV.scala 172:21]
    end
    if (reset) begin // @[Cordic_LV.scala 161:38]
      y_flag_reg_7 <= 1'h0; // @[Cordic_LV.scala 161:38]
    end else begin
      y_flag_reg_7 <= y_flag_reg_6; // @[Cordic_LV.scala 172:21]
    end
    if (reset) begin // @[Cordic_LV.scala 161:38]
      y_flag_reg_8 <= 1'h0; // @[Cordic_LV.scala 161:38]
    end else begin
      y_flag_reg_8 <= y_flag_reg_7; // @[Cordic_LV.scala 172:21]
    end
    if (reset) begin // @[Cordic_LV.scala 161:38]
      y_flag_reg_9 <= 1'h0; // @[Cordic_LV.scala 161:38]
    end else begin
      y_flag_reg_9 <= y_flag_reg_8; // @[Cordic_LV.scala 172:21]
    end
    if (reset) begin // @[Cordic_LV.scala 161:38]
      y_flag_reg_10 <= 1'h0; // @[Cordic_LV.scala 161:38]
    end else begin
      y_flag_reg_10 <= y_flag_reg_9; // @[Cordic_LV.scala 172:21]
    end
    if (reset) begin // @[Cordic_LV.scala 161:38]
      y_flag_reg_11 <= 1'h0; // @[Cordic_LV.scala 161:38]
    end else begin
      y_flag_reg_11 <= y_flag_reg_10; // @[Cordic_LV.scala 172:21]
    end
    if (reset) begin // @[Cordic_LV.scala 161:38]
      y_flag_reg_12 <= 1'h0; // @[Cordic_LV.scala 161:38]
    end else begin
      y_flag_reg_12 <= y_flag_reg_11; // @[Cordic_LV.scala 172:21]
    end
    if (reset) begin // @[Cordic_LV.scala 161:38]
      y_flag_reg_13 <= 1'h0; // @[Cordic_LV.scala 161:38]
    end else begin
      y_flag_reg_13 <= y_flag_reg_12; // @[Cordic_LV.scala 172:21]
    end
    if (reset) begin // @[Cordic_LV.scala 161:38]
      y_flag_reg_14 <= 1'h0; // @[Cordic_LV.scala 161:38]
    end else begin
      y_flag_reg_14 <= y_flag_reg_13; // @[Cordic_LV.scala 172:21]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  x_cnt_reg_0 = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  x_cnt_reg_1 = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  x_cnt_reg_2 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  x_cnt_reg_3 = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  x_cnt_reg_4 = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  x_cnt_reg_5 = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  x_cnt_reg_6 = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  x_cnt_reg_7 = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  x_cnt_reg_8 = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  x_cnt_reg_9 = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
  x_cnt_reg_10 = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  x_cnt_reg_11 = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  x_cnt_reg_12 = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  x_cnt_reg_13 = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  x_cnt_reg_14 = _RAND_14[5:0];
  _RAND_15 = {1{`RANDOM}};
  x_flag_reg_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  x_flag_reg_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  x_flag_reg_2 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  x_flag_reg_3 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  x_flag_reg_4 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  x_flag_reg_5 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  x_flag_reg_6 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  x_flag_reg_7 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  x_flag_reg_8 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  x_flag_reg_9 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  x_flag_reg_10 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  x_flag_reg_11 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  x_flag_reg_12 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  x_flag_reg_13 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  x_flag_reg_14 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  y_cnt_reg_0 = _RAND_30[5:0];
  _RAND_31 = {1{`RANDOM}};
  y_cnt_reg_1 = _RAND_31[5:0];
  _RAND_32 = {1{`RANDOM}};
  y_cnt_reg_2 = _RAND_32[5:0];
  _RAND_33 = {1{`RANDOM}};
  y_cnt_reg_3 = _RAND_33[5:0];
  _RAND_34 = {1{`RANDOM}};
  y_cnt_reg_4 = _RAND_34[5:0];
  _RAND_35 = {1{`RANDOM}};
  y_cnt_reg_5 = _RAND_35[5:0];
  _RAND_36 = {1{`RANDOM}};
  y_cnt_reg_6 = _RAND_36[5:0];
  _RAND_37 = {1{`RANDOM}};
  y_cnt_reg_7 = _RAND_37[5:0];
  _RAND_38 = {1{`RANDOM}};
  y_cnt_reg_8 = _RAND_38[5:0];
  _RAND_39 = {1{`RANDOM}};
  y_cnt_reg_9 = _RAND_39[5:0];
  _RAND_40 = {1{`RANDOM}};
  y_cnt_reg_10 = _RAND_40[5:0];
  _RAND_41 = {1{`RANDOM}};
  y_cnt_reg_11 = _RAND_41[5:0];
  _RAND_42 = {1{`RANDOM}};
  y_cnt_reg_12 = _RAND_42[5:0];
  _RAND_43 = {1{`RANDOM}};
  y_cnt_reg_13 = _RAND_43[5:0];
  _RAND_44 = {1{`RANDOM}};
  y_cnt_reg_14 = _RAND_44[5:0];
  _RAND_45 = {1{`RANDOM}};
  y_flag_reg_0 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  y_flag_reg_1 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  y_flag_reg_2 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  y_flag_reg_3 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  y_flag_reg_4 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  y_flag_reg_5 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  y_flag_reg_6 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  y_flag_reg_7 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  y_flag_reg_8 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  y_flag_reg_9 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  y_flag_reg_10 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  y_flag_reg_11 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  y_flag_reg_12 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  y_flag_reg_13 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  y_flag_reg_14 = _RAND_59[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cordic_sin_cos_expand(
  input         clock,
  input         reset,
  input  [63:0] io_theta,
  output [63:0] io_sin,
  output [63:0] io_cos
);
  wire  cordic_unit_clock; // @[Cordic_CR.scala 171:29]
  wire  cordic_unit_reset; // @[Cordic_CR.scala 171:29]
  wire [63:0] cordic_unit_io_theta; // @[Cordic_CR.scala 171:29]
  wire [63:0] cordic_unit_io_sin; // @[Cordic_CR.scala 171:29]
  wire [63:0] cordic_unit_io_cos; // @[Cordic_CR.scala 171:29]
  wire [63:0] _T_3 = $signed(io_theta) + 64'sh16800000000; // @[Cordic_CR.scala 230:21]
  wire  index__0 = $signed(_T_3) < -64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 230:72 231:18 233:18]
  wire [63:0] _T_7 = $signed(io_theta) + 64'sh2d000000000; // @[Cordic_CR.scala 230:21]
  wire  index__1 = $signed(_T_7) < -64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 230:72 231:18 233:18]
  wire [63:0] _T_11 = $signed(io_theta) + 64'sh43800000000; // @[Cordic_CR.scala 230:21]
  wire  index__2 = $signed(_T_11) < -64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 230:72 231:18 233:18]
  wire [63:0] _T_15 = $signed(io_theta) + 64'sh5a000000000; // @[Cordic_CR.scala 230:21]
  wire  index__3 = $signed(_T_15) < -64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 230:72 231:18 233:18]
  wire [63:0] _T_19 = $signed(io_theta) + 64'sh70800000000; // @[Cordic_CR.scala 230:21]
  wire  index__4 = $signed(_T_19) < -64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 230:72 231:18 233:18]
  wire [63:0] _T_23 = $signed(io_theta) + 64'sh87000000000; // @[Cordic_CR.scala 230:21]
  wire  index__5 = $signed(_T_23) < -64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 230:72 231:18 233:18]
  wire [63:0] _T_27 = $signed(io_theta) + 64'sh9d800000000; // @[Cordic_CR.scala 230:21]
  wire  index__6 = $signed(_T_27) < -64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 230:72 231:18 233:18]
  wire [63:0] _T_31 = $signed(io_theta) + 64'shb4000000000; // @[Cordic_CR.scala 230:21]
  wire  index__7 = $signed(_T_31) < -64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 230:72 231:18 233:18]
  wire [63:0] _T_35 = $signed(io_theta) + 64'shca800000000; // @[Cordic_CR.scala 230:21]
  wire  index__8 = $signed(_T_35) < -64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 230:72 231:18 233:18]
  wire [63:0] _T_39 = $signed(io_theta) + 64'she1000000000; // @[Cordic_CR.scala 230:21]
  wire  index__9 = $signed(_T_39) < -64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 230:72 231:18 233:18]
  wire [9:0] _temp_cnt_T = {index__9,index__8,index__7,index__6,index__5,index__4,index__3,index__2,index__1,index__0}; // @[Cordic_CR.scala 237:48]
  wire [3:0] _temp_cnt_T_11 = _temp_cnt_T[8] ? 4'h8 : 4'h9; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_12 = _temp_cnt_T[7] ? 4'h7 : _temp_cnt_T_11; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_13 = _temp_cnt_T[6] ? 4'h6 : _temp_cnt_T_12; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_14 = _temp_cnt_T[5] ? 4'h5 : _temp_cnt_T_13; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_15 = _temp_cnt_T[4] ? 4'h4 : _temp_cnt_T_14; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_16 = _temp_cnt_T[3] ? 4'h3 : _temp_cnt_T_15; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_17 = _temp_cnt_T[2] ? 4'h2 : _temp_cnt_T_16; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_18 = _temp_cnt_T[1] ? 4'h1 : _temp_cnt_T_17; // @[Mux.scala 47:70]
  wire [3:0] temp_cnt = _temp_cnt_T[0] ? 4'h0 : _temp_cnt_T_18; // @[Mux.scala 47:70]
  wire [63:0] _GEN_11 = 4'h1 == temp_cnt ? $signed(64'sh2d000000000) : $signed(64'sh16800000000); // @[Cordic_CR.scala 238:{28,28}]
  wire [63:0] _GEN_12 = 4'h2 == temp_cnt ? $signed(64'sh43800000000) : $signed(_GEN_11); // @[Cordic_CR.scala 238:{28,28}]
  wire [63:0] _GEN_13 = 4'h3 == temp_cnt ? $signed(64'sh5a000000000) : $signed(_GEN_12); // @[Cordic_CR.scala 238:{28,28}]
  wire [63:0] _GEN_14 = 4'h4 == temp_cnt ? $signed(64'sh70800000000) : $signed(_GEN_13); // @[Cordic_CR.scala 238:{28,28}]
  wire [63:0] _GEN_15 = 4'h5 == temp_cnt ? $signed(64'sh87000000000) : $signed(_GEN_14); // @[Cordic_CR.scala 238:{28,28}]
  wire [63:0] _GEN_16 = 4'h6 == temp_cnt ? $signed(64'sh9d800000000) : $signed(_GEN_15); // @[Cordic_CR.scala 238:{28,28}]
  wire [63:0] _GEN_17 = 4'h7 == temp_cnt ? $signed(64'shb4000000000) : $signed(_GEN_16); // @[Cordic_CR.scala 238:{28,28}]
  wire [63:0] _GEN_18 = 4'h8 == temp_cnt ? $signed(64'shca800000000) : $signed(_GEN_17); // @[Cordic_CR.scala 238:{28,28}]
  wire [63:0] _GEN_19 = 4'h9 == temp_cnt ? $signed(64'she1000000000) : $signed(_GEN_18); // @[Cordic_CR.scala 238:{28,28}]
  wire [63:0] _real_theta_T_2 = $signed(io_theta) + $signed(_GEN_19); // @[Cordic_CR.scala 238:28]
  wire [63:0] _T_44 = $signed(io_theta) - 64'sh16800000000; // @[Cordic_CR.scala 243:21]
  wire  index_1_0 = $signed(_T_44) > 64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 243:71 244:18 246:18]
  wire [63:0] _T_48 = $signed(io_theta) - 64'sh2d000000000; // @[Cordic_CR.scala 243:21]
  wire  index_1_1 = $signed(_T_48) > 64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 243:71 244:18 246:18]
  wire [63:0] _T_52 = $signed(io_theta) - 64'sh43800000000; // @[Cordic_CR.scala 243:21]
  wire  index_1_2 = $signed(_T_52) > 64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 243:71 244:18 246:18]
  wire [63:0] _T_56 = $signed(io_theta) - 64'sh5a000000000; // @[Cordic_CR.scala 243:21]
  wire  index_1_3 = $signed(_T_56) > 64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 243:71 244:18 246:18]
  wire [63:0] _T_60 = $signed(io_theta) - 64'sh70800000000; // @[Cordic_CR.scala 243:21]
  wire  index_1_4 = $signed(_T_60) > 64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 243:71 244:18 246:18]
  wire [63:0] _T_64 = $signed(io_theta) - 64'sh87000000000; // @[Cordic_CR.scala 243:21]
  wire  index_1_5 = $signed(_T_64) > 64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 243:71 244:18 246:18]
  wire [63:0] _T_68 = $signed(io_theta) - 64'sh9d800000000; // @[Cordic_CR.scala 243:21]
  wire  index_1_6 = $signed(_T_68) > 64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 243:71 244:18 246:18]
  wire [63:0] _T_72 = $signed(io_theta) - 64'shb4000000000; // @[Cordic_CR.scala 243:21]
  wire  index_1_7 = $signed(_T_72) > 64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 243:71 244:18 246:18]
  wire [63:0] _T_76 = $signed(io_theta) - 64'shca800000000; // @[Cordic_CR.scala 243:21]
  wire  index_1_8 = $signed(_T_76) > 64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 243:71 244:18 246:18]
  wire [63:0] _T_80 = $signed(io_theta) - 64'she1000000000; // @[Cordic_CR.scala 243:21]
  wire  index_1_9 = $signed(_T_80) > 64'sh16800000000 ? 1'h0 : 1'h1; // @[Cordic_CR.scala 243:71 244:18 246:18]
  wire [9:0] _temp_cnt_T_19 = {index_1_9,index_1_8,index_1_7,index_1_6,index_1_5,index_1_4,index_1_3,index_1_2,index_1_1
    ,index_1_0}; // @[Cordic_CR.scala 250:48]
  wire [3:0] _temp_cnt_T_30 = _temp_cnt_T_19[8] ? 4'h8 : 4'h9; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_31 = _temp_cnt_T_19[7] ? 4'h7 : _temp_cnt_T_30; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_32 = _temp_cnt_T_19[6] ? 4'h6 : _temp_cnt_T_31; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_33 = _temp_cnt_T_19[5] ? 4'h5 : _temp_cnt_T_32; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_34 = _temp_cnt_T_19[4] ? 4'h4 : _temp_cnt_T_33; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_35 = _temp_cnt_T_19[3] ? 4'h3 : _temp_cnt_T_34; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_36 = _temp_cnt_T_19[2] ? 4'h2 : _temp_cnt_T_35; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_37 = _temp_cnt_T_19[1] ? 4'h1 : _temp_cnt_T_36; // @[Mux.scala 47:70]
  wire [3:0] temp_cnt_1 = _temp_cnt_T_19[0] ? 4'h0 : _temp_cnt_T_37; // @[Mux.scala 47:70]
  wire [63:0] _GEN_31 = 4'h1 == temp_cnt_1 ? $signed(64'sh2d000000000) : $signed(64'sh16800000000); // @[Cordic_CR.scala 251:{28,28}]
  wire [63:0] _GEN_32 = 4'h2 == temp_cnt_1 ? $signed(64'sh43800000000) : $signed(_GEN_31); // @[Cordic_CR.scala 251:{28,28}]
  wire [63:0] _GEN_33 = 4'h3 == temp_cnt_1 ? $signed(64'sh5a000000000) : $signed(_GEN_32); // @[Cordic_CR.scala 251:{28,28}]
  wire [63:0] _GEN_34 = 4'h4 == temp_cnt_1 ? $signed(64'sh70800000000) : $signed(_GEN_33); // @[Cordic_CR.scala 251:{28,28}]
  wire [63:0] _GEN_35 = 4'h5 == temp_cnt_1 ? $signed(64'sh87000000000) : $signed(_GEN_34); // @[Cordic_CR.scala 251:{28,28}]
  wire [63:0] _GEN_36 = 4'h6 == temp_cnt_1 ? $signed(64'sh9d800000000) : $signed(_GEN_35); // @[Cordic_CR.scala 251:{28,28}]
  wire [63:0] _GEN_37 = 4'h7 == temp_cnt_1 ? $signed(64'shb4000000000) : $signed(_GEN_36); // @[Cordic_CR.scala 251:{28,28}]
  wire [63:0] _GEN_38 = 4'h8 == temp_cnt_1 ? $signed(64'shca800000000) : $signed(_GEN_37); // @[Cordic_CR.scala 251:{28,28}]
  wire [63:0] _GEN_39 = 4'h9 == temp_cnt_1 ? $signed(64'she1000000000) : $signed(_GEN_38); // @[Cordic_CR.scala 251:{28,28}]
  wire [63:0] _real_theta_T_5 = $signed(io_theta) - $signed(_GEN_39); // @[Cordic_CR.scala 251:28]
  wire [63:0] _GEN_40 = $signed(io_theta) > 64'sh16800000000 ? $signed(_real_theta_T_5) : $signed(io_theta); // @[Cordic_CR.scala 239:82 251:16 253:16]
  cordic_sin_cos cordic_unit ( // @[Cordic_CR.scala 171:29]
    .clock(cordic_unit_clock),
    .reset(cordic_unit_reset),
    .io_theta(cordic_unit_io_theta),
    .io_sin(cordic_unit_io_sin),
    .io_cos(cordic_unit_io_cos)
  );
  assign io_sin = cordic_unit_io_sin; // @[Cordic_CR.scala 256:10]
  assign io_cos = cordic_unit_io_cos; // @[Cordic_CR.scala 257:10]
  assign cordic_unit_clock = clock;
  assign cordic_unit_reset = reset;
  assign cordic_unit_io_theta = $signed(io_theta) < -64'sh16800000000 ? $signed(_real_theta_T_2) : $signed(_GEN_40); // @[Cordic_CR.scala 226:77 238:16]
endmodule
module ComplexMul(
  input  [63:0] io_op1_re,
  input  [63:0] io_op1_im,
  input  [63:0] io_op2_re,
  input  [63:0] io_op2_im,
  output [63:0] io_res_re,
  output [63:0] io_res_im
);
  wire [63:0] _k1_T_2 = $signed(io_op1_re) + $signed(io_op1_im); // @[Complex_Operater.scala 38:35]
  wire [127:0] k1 = $signed(io_op2_re) * $signed(_k1_T_2); // @[Complex_Operater.scala 38:22]
  wire [63:0] _k2_T_2 = $signed(io_op2_im) - $signed(io_op2_re); // @[Complex_Operater.scala 39:35]
  wire [127:0] k2 = $signed(io_op1_re) * $signed(_k2_T_2); // @[Complex_Operater.scala 39:22]
  wire [63:0] _k3_T_2 = $signed(io_op2_re) + $signed(io_op2_im); // @[Complex_Operater.scala 40:35]
  wire [127:0] k3 = $signed(io_op1_im) * $signed(_k3_T_2); // @[Complex_Operater.scala 40:22]
  wire [127:0] _io_res_re_T_2 = $signed(k1) - $signed(k3); // @[Complex_Operater.scala 41:19]
  wire [127:0] _io_res_im_T_2 = $signed(k1) + $signed(k2); // @[Complex_Operater.scala 42:19]
  wire [95:0] _GEN_0 = _io_res_re_T_2[127:32]; // @[Complex_Operater.scala 41:13]
  wire [95:0] _GEN_2 = _io_res_im_T_2[127:32]; // @[Complex_Operater.scala 42:13]
  assign io_res_re = _GEN_0[63:0]; // @[Complex_Operater.scala 41:13]
  assign io_res_im = _GEN_2[63:0]; // @[Complex_Operater.scala 42:13]
endmodule
module matrix_vlaue_mul(
  input  [63:0] io_matrixIn_1_re,
  input  [63:0] io_matrixIn_1_im,
  input  [63:0] io_valueIn_re,
  input  [63:0] io_valueIn_im,
  output [63:0] io_matrixOut_0_re,
  output [63:0] io_matrixOut_0_im,
  output [63:0] io_matrixOut_1_re,
  output [63:0] io_matrixOut_1_im
);
  wire [63:0] io_matrixOut_0_mul_io_op1_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_0_mul_io_op1_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_0_mul_io_op2_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_0_mul_io_op2_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_0_mul_io_res_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_0_mul_io_res_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_1_mul_io_op1_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_1_mul_io_op1_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_1_mul_io_op2_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_1_mul_io_op2_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_1_mul_io_res_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_1_mul_io_res_im; // @[Complex_Operater.scala 47:21]
  ComplexMul io_matrixOut_0_mul ( // @[Complex_Operater.scala 47:21]
    .io_op1_re(io_matrixOut_0_mul_io_op1_re),
    .io_op1_im(io_matrixOut_0_mul_io_op1_im),
    .io_op2_re(io_matrixOut_0_mul_io_op2_re),
    .io_op2_im(io_matrixOut_0_mul_io_op2_im),
    .io_res_re(io_matrixOut_0_mul_io_res_re),
    .io_res_im(io_matrixOut_0_mul_io_res_im)
  );
  ComplexMul io_matrixOut_1_mul ( // @[Complex_Operater.scala 47:21]
    .io_op1_re(io_matrixOut_1_mul_io_op1_re),
    .io_op1_im(io_matrixOut_1_mul_io_op1_im),
    .io_op2_re(io_matrixOut_1_mul_io_op2_re),
    .io_op2_im(io_matrixOut_1_mul_io_op2_im),
    .io_res_re(io_matrixOut_1_mul_io_res_re),
    .io_res_im(io_matrixOut_1_mul_io_res_im)
  );
  assign io_matrixOut_0_re = io_matrixOut_0_mul_io_res_re; // @[Kronecker_V1.scala 24:21]
  assign io_matrixOut_0_im = io_matrixOut_0_mul_io_res_im; // @[Kronecker_V1.scala 24:21]
  assign io_matrixOut_1_re = io_matrixOut_1_mul_io_res_re; // @[Kronecker_V1.scala 24:21]
  assign io_matrixOut_1_im = io_matrixOut_1_mul_io_res_im; // @[Kronecker_V1.scala 24:21]
  assign io_matrixOut_0_mul_io_op1_re = 64'sh100000000; // @[Complex_Operater.scala 48:16]
  assign io_matrixOut_0_mul_io_op1_im = 64'sh0; // @[Complex_Operater.scala 48:16]
  assign io_matrixOut_0_mul_io_op2_re = io_valueIn_re; // @[Complex_Operater.scala 49:16]
  assign io_matrixOut_0_mul_io_op2_im = io_valueIn_im; // @[Complex_Operater.scala 49:16]
  assign io_matrixOut_1_mul_io_op1_re = io_matrixIn_1_re; // @[Complex_Operater.scala 48:16]
  assign io_matrixOut_1_mul_io_op1_im = io_matrixIn_1_im; // @[Complex_Operater.scala 48:16]
  assign io_matrixOut_1_mul_io_op2_re = io_valueIn_re; // @[Complex_Operater.scala 49:16]
  assign io_matrixOut_1_mul_io_op2_im = io_valueIn_im; // @[Complex_Operater.scala 49:16]
endmodule
module kronecker_v1(
  input  [63:0] io_matrixA_1_re,
  input  [63:0] io_matrixA_1_im,
  input  [63:0] io_matrixB_1_re,
  input  [63:0] io_matrixB_1_im,
  output [63:0] io_matrixOut_0_re,
  output [63:0] io_matrixOut_0_im,
  output [63:0] io_matrixOut_1_re,
  output [63:0] io_matrixOut_1_im,
  output [63:0] io_matrixOut_2_re,
  output [63:0] io_matrixOut_2_im,
  output [63:0] io_matrixOut_3_re,
  output [63:0] io_matrixOut_3_im
);
  wire [63:0] unit_io_matrixIn_1_re; // @[Kronecker_V1.scala 39:22]
  wire [63:0] unit_io_matrixIn_1_im; // @[Kronecker_V1.scala 39:22]
  wire [63:0] unit_io_valueIn_re; // @[Kronecker_V1.scala 39:22]
  wire [63:0] unit_io_valueIn_im; // @[Kronecker_V1.scala 39:22]
  wire [63:0] unit_io_matrixOut_0_re; // @[Kronecker_V1.scala 39:22]
  wire [63:0] unit_io_matrixOut_0_im; // @[Kronecker_V1.scala 39:22]
  wire [63:0] unit_io_matrixOut_1_re; // @[Kronecker_V1.scala 39:22]
  wire [63:0] unit_io_matrixOut_1_im; // @[Kronecker_V1.scala 39:22]
  wire [63:0] unit_1_io_matrixIn_1_re; // @[Kronecker_V1.scala 39:22]
  wire [63:0] unit_1_io_matrixIn_1_im; // @[Kronecker_V1.scala 39:22]
  wire [63:0] unit_1_io_valueIn_re; // @[Kronecker_V1.scala 39:22]
  wire [63:0] unit_1_io_valueIn_im; // @[Kronecker_V1.scala 39:22]
  wire [63:0] unit_1_io_matrixOut_0_re; // @[Kronecker_V1.scala 39:22]
  wire [63:0] unit_1_io_matrixOut_0_im; // @[Kronecker_V1.scala 39:22]
  wire [63:0] unit_1_io_matrixOut_1_re; // @[Kronecker_V1.scala 39:22]
  wire [63:0] unit_1_io_matrixOut_1_im; // @[Kronecker_V1.scala 39:22]
  matrix_vlaue_mul unit ( // @[Kronecker_V1.scala 39:22]
    .io_matrixIn_1_re(unit_io_matrixIn_1_re),
    .io_matrixIn_1_im(unit_io_matrixIn_1_im),
    .io_valueIn_re(unit_io_valueIn_re),
    .io_valueIn_im(unit_io_valueIn_im),
    .io_matrixOut_0_re(unit_io_matrixOut_0_re),
    .io_matrixOut_0_im(unit_io_matrixOut_0_im),
    .io_matrixOut_1_re(unit_io_matrixOut_1_re),
    .io_matrixOut_1_im(unit_io_matrixOut_1_im)
  );
  matrix_vlaue_mul unit_1 ( // @[Kronecker_V1.scala 39:22]
    .io_matrixIn_1_re(unit_1_io_matrixIn_1_re),
    .io_matrixIn_1_im(unit_1_io_matrixIn_1_im),
    .io_valueIn_re(unit_1_io_valueIn_re),
    .io_valueIn_im(unit_1_io_valueIn_im),
    .io_matrixOut_0_re(unit_1_io_matrixOut_0_re),
    .io_matrixOut_0_im(unit_1_io_matrixOut_0_im),
    .io_matrixOut_1_re(unit_1_io_matrixOut_1_re),
    .io_matrixOut_1_im(unit_1_io_matrixOut_1_im)
  );
  assign io_matrixOut_0_re = unit_io_matrixOut_0_re; // @[Kronecker_V1.scala 67:29 68:19]
  assign io_matrixOut_0_im = unit_io_matrixOut_0_im; // @[Kronecker_V1.scala 67:29 68:19]
  assign io_matrixOut_1_re = unit_io_matrixOut_1_re; // @[Kronecker_V1.scala 67:29 68:19]
  assign io_matrixOut_1_im = unit_io_matrixOut_1_im; // @[Kronecker_V1.scala 67:29 68:19]
  assign io_matrixOut_2_re = unit_1_io_matrixOut_0_re; // @[Kronecker_V1.scala 67:29 68:19]
  assign io_matrixOut_2_im = unit_1_io_matrixOut_0_im; // @[Kronecker_V1.scala 67:29 68:19]
  assign io_matrixOut_3_re = unit_1_io_matrixOut_1_re; // @[Kronecker_V1.scala 67:29 68:19]
  assign io_matrixOut_3_im = unit_1_io_matrixOut_1_im; // @[Kronecker_V1.scala 67:29 68:19]
  assign unit_io_matrixIn_1_re = io_matrixB_1_re; // @[Kronecker_V1.scala 40:22]
  assign unit_io_matrixIn_1_im = io_matrixB_1_im; // @[Kronecker_V1.scala 40:22]
  assign unit_io_valueIn_re = 64'sh100000000; // @[Kronecker_V1.scala 41:21]
  assign unit_io_valueIn_im = 64'sh0; // @[Kronecker_V1.scala 41:21]
  assign unit_1_io_matrixIn_1_re = io_matrixB_1_re; // @[Kronecker_V1.scala 40:22]
  assign unit_1_io_matrixIn_1_im = io_matrixB_1_im; // @[Kronecker_V1.scala 40:22]
  assign unit_1_io_valueIn_re = io_matrixA_1_re; // @[Kronecker_V1.scala 41:21]
  assign unit_1_io_valueIn_im = io_matrixA_1_im; // @[Kronecker_V1.scala 41:21]
endmodule
module space_time_steering_vector(
  input         clock,
  input         reset,
  input  [63:0] io_theta,
  input  [63:0] io_psi,
  input  [63:0] io_d,
  input  [63:0] io_lambda,
  input  [63:0] io_v,
  input  [63:0] io_T,
  output [63:0] io_matrixOut_0_re,
  output [63:0] io_matrixOut_0_im,
  output [63:0] io_matrixOut_1_re,
  output [63:0] io_matrixOut_1_im,
  output [63:0] io_matrixOut_2_re,
  output [63:0] io_matrixOut_2_im,
  output [63:0] io_matrixOut_3_re,
  output [63:0] io_matrixOut_3_im
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
`endif // RANDOMIZE_REG_INIT
  wire  cordic_unit_clock; // @[Cordic_CR.scala 171:29]
  wire  cordic_unit_reset; // @[Cordic_CR.scala 171:29]
  wire [63:0] cordic_unit_io_theta; // @[Cordic_CR.scala 171:29]
  wire [63:0] cordic_unit_io_sin; // @[Cordic_CR.scala 171:29]
  wire [63:0] cordic_unit_io_cos; // @[Cordic_CR.scala 171:29]
  wire  cordic_unit_1_clock; // @[Cordic_CR.scala 171:29]
  wire  cordic_unit_1_reset; // @[Cordic_CR.scala 171:29]
  wire [63:0] cordic_unit_1_io_theta; // @[Cordic_CR.scala 171:29]
  wire [63:0] cordic_unit_1_io_sin; // @[Cordic_CR.scala 171:29]
  wire [63:0] cordic_unit_1_io_cos; // @[Cordic_CR.scala 171:29]
  wire  lambda_divide_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  lambda_divide_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] lambda_divide_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] lambda_divide_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] lambda_divide_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  cordic_unit_2_clock; // @[Cordic_CR.scala 271:29]
  wire  cordic_unit_2_reset; // @[Cordic_CR.scala 271:29]
  wire [63:0] cordic_unit_2_io_theta; // @[Cordic_CR.scala 271:29]
  wire [63:0] cordic_unit_2_io_sin; // @[Cordic_CR.scala 271:29]
  wire [63:0] cordic_unit_2_io_cos; // @[Cordic_CR.scala 271:29]
  wire  cordic_unit_3_clock; // @[Cordic_CR.scala 271:29]
  wire  cordic_unit_3_reset; // @[Cordic_CR.scala 271:29]
  wire [63:0] cordic_unit_3_io_theta; // @[Cordic_CR.scala 271:29]
  wire [63:0] cordic_unit_3_io_sin; // @[Cordic_CR.scala 271:29]
  wire [63:0] cordic_unit_3_io_cos; // @[Cordic_CR.scala 271:29]
  wire [63:0] unit_io_matrixA_1_re; // @[Kronecker_V1.scala 92:22]
  wire [63:0] unit_io_matrixA_1_im; // @[Kronecker_V1.scala 92:22]
  wire [63:0] unit_io_matrixB_1_re; // @[Kronecker_V1.scala 92:22]
  wire [63:0] unit_io_matrixB_1_im; // @[Kronecker_V1.scala 92:22]
  wire [63:0] unit_io_matrixOut_0_re; // @[Kronecker_V1.scala 92:22]
  wire [63:0] unit_io_matrixOut_0_im; // @[Kronecker_V1.scala 92:22]
  wire [63:0] unit_io_matrixOut_1_re; // @[Kronecker_V1.scala 92:22]
  wire [63:0] unit_io_matrixOut_1_im; // @[Kronecker_V1.scala 92:22]
  wire [63:0] unit_io_matrixOut_2_re; // @[Kronecker_V1.scala 92:22]
  wire [63:0] unit_io_matrixOut_2_im; // @[Kronecker_V1.scala 92:22]
  wire [63:0] unit_io_matrixOut_3_re; // @[Kronecker_V1.scala 92:22]
  wire [63:0] unit_io_matrixOut_3_im; // @[Kronecker_V1.scala 92:22]
  reg [63:0] reg_d_0; // @[Space_Time_Steering_Vector.scala 40:39]
  reg [63:0] reg_d_1; // @[Space_Time_Steering_Vector.scala 40:39]
  reg [63:0] reg_d_2; // @[Space_Time_Steering_Vector.scala 40:39]
  reg [63:0] reg_d_3; // @[Space_Time_Steering_Vector.scala 40:39]
  reg [63:0] reg_d_4; // @[Space_Time_Steering_Vector.scala 40:39]
  reg [63:0] reg_d_5; // @[Space_Time_Steering_Vector.scala 40:39]
  reg [63:0] reg_d_6; // @[Space_Time_Steering_Vector.scala 40:39]
  reg [63:0] reg_d_7; // @[Space_Time_Steering_Vector.scala 40:39]
  reg [63:0] reg_d_8; // @[Space_Time_Steering_Vector.scala 40:39]
  reg [63:0] reg_d_9; // @[Space_Time_Steering_Vector.scala 40:39]
  reg [63:0] reg_d_10; // @[Space_Time_Steering_Vector.scala 40:39]
  reg [63:0] reg_d_11; // @[Space_Time_Steering_Vector.scala 40:39]
  reg [63:0] reg_d_12; // @[Space_Time_Steering_Vector.scala 40:39]
  reg [63:0] reg_d_13; // @[Space_Time_Steering_Vector.scala 40:39]
  reg [63:0] reg_d_14; // @[Space_Time_Steering_Vector.scala 40:39]
  reg [63:0] reg_v_0; // @[Space_Time_Steering_Vector.scala 41:39]
  reg [63:0] reg_v_1; // @[Space_Time_Steering_Vector.scala 41:39]
  reg [63:0] reg_v_2; // @[Space_Time_Steering_Vector.scala 41:39]
  reg [63:0] reg_v_3; // @[Space_Time_Steering_Vector.scala 41:39]
  reg [63:0] reg_v_4; // @[Space_Time_Steering_Vector.scala 41:39]
  reg [63:0] reg_v_5; // @[Space_Time_Steering_Vector.scala 41:39]
  reg [63:0] reg_v_6; // @[Space_Time_Steering_Vector.scala 41:39]
  reg [63:0] reg_v_7; // @[Space_Time_Steering_Vector.scala 41:39]
  reg [63:0] reg_v_8; // @[Space_Time_Steering_Vector.scala 41:39]
  reg [63:0] reg_v_9; // @[Space_Time_Steering_Vector.scala 41:39]
  reg [63:0] reg_v_10; // @[Space_Time_Steering_Vector.scala 41:39]
  reg [63:0] reg_v_11; // @[Space_Time_Steering_Vector.scala 41:39]
  reg [63:0] reg_v_12; // @[Space_Time_Steering_Vector.scala 41:39]
  reg [63:0] reg_v_13; // @[Space_Time_Steering_Vector.scala 41:39]
  reg [63:0] reg_v_14; // @[Space_Time_Steering_Vector.scala 41:39]
  reg [63:0] reg_T_0; // @[Space_Time_Steering_Vector.scala 42:39]
  reg [63:0] reg_T_1; // @[Space_Time_Steering_Vector.scala 42:39]
  reg [63:0] reg_T_2; // @[Space_Time_Steering_Vector.scala 42:39]
  reg [63:0] reg_T_3; // @[Space_Time_Steering_Vector.scala 42:39]
  reg [63:0] reg_T_4; // @[Space_Time_Steering_Vector.scala 42:39]
  reg [63:0] reg_T_5; // @[Space_Time_Steering_Vector.scala 42:39]
  reg [63:0] reg_T_6; // @[Space_Time_Steering_Vector.scala 42:39]
  reg [63:0] reg_T_7; // @[Space_Time_Steering_Vector.scala 42:39]
  reg [63:0] reg_T_8; // @[Space_Time_Steering_Vector.scala 42:39]
  reg [63:0] reg_T_9; // @[Space_Time_Steering_Vector.scala 42:39]
  reg [63:0] reg_T_10; // @[Space_Time_Steering_Vector.scala 42:39]
  reg [63:0] reg_T_11; // @[Space_Time_Steering_Vector.scala 42:39]
  reg [63:0] reg_T_12; // @[Space_Time_Steering_Vector.scala 42:39]
  reg [63:0] reg_T_13; // @[Space_Time_Steering_Vector.scala 42:39]
  reg [63:0] reg_T_14; // @[Space_Time_Steering_Vector.scala 42:39]
  wire [127:0] _fs_T = $signed(reg_d_14) * $signed(cordic_unit_io_cos); // @[Space_Time_Steering_Vector.scala 61:50]
  wire [191:0] _fs_T_1 = $signed(_fs_T) * $signed(cordic_unit_1_io_cos); // @[Space_Time_Steering_Vector.scala 61:62]
  wire [255:0] fs = $signed(_fs_T_1) * $signed(lambda_divide_divide_io_z); // @[Space_Time_Steering_Vector.scala 61:72]
  wire [127:0] _fd_T = $signed(reg_v_14) * $signed(reg_T_14); // @[Space_Time_Steering_Vector.scala 62:51]
  wire [191:0] _fd_T_1 = $signed(_fd_T) * $signed(cordic_unit_io_cos); // @[Space_Time_Steering_Vector.scala 62:79]
  wire [255:0] _fd_T_2 = $signed(_fd_T_1) * $signed(cordic_unit_1_io_cos); // @[Space_Time_Steering_Vector.scala 62:91]
  wire [319:0] _fd_T_3 = $signed(_fd_T_2) * $signed(lambda_divide_divide_io_z); // @[Space_Time_Steering_Vector.scala 62:101]
  wire [320:0] fd = {$signed(_fd_T_3), 1'h0}; // @[Space_Time_Steering_Vector.scala 62:118]
  wire [319:0] cal_in = 64'sh16800000000 * $signed(fs); // @[Space_Time_Steering_Vector.scala 74:103]
  wire [384:0] cal_in_1 = 64'sh16800000000 * $signed(fd); // @[Space_Time_Steering_Vector.scala 81:103]
  wire [191:0] _GEN_4 = cal_in[319:128]; // @[Cordic_CR.scala 272:26]
  wire [224:0] _GEN_6 = cal_in_1[384:160]; // @[Cordic_CR.scala 272:26]
  cordic_sin_cos cordic_unit ( // @[Cordic_CR.scala 171:29]
    .clock(cordic_unit_clock),
    .reset(cordic_unit_reset),
    .io_theta(cordic_unit_io_theta),
    .io_sin(cordic_unit_io_sin),
    .io_cos(cordic_unit_io_cos)
  );
  cordic_sin_cos cordic_unit_1 ( // @[Cordic_CR.scala 171:29]
    .clock(cordic_unit_1_clock),
    .reset(cordic_unit_1_reset),
    .io_theta(cordic_unit_1_io_theta),
    .io_sin(cordic_unit_1_io_sin),
    .io_cos(cordic_unit_1_io_cos)
  );
  cordic_divide lambda_divide_divide ( // @[Cordic_LV.scala 211:24]
    .clock(lambda_divide_divide_clock),
    .reset(lambda_divide_divide_reset),
    .io_x(lambda_divide_divide_io_x),
    .io_y(lambda_divide_divide_io_y),
    .io_z(lambda_divide_divide_io_z)
  );
  cordic_sin_cos_expand cordic_unit_2 ( // @[Cordic_CR.scala 271:29]
    .clock(cordic_unit_2_clock),
    .reset(cordic_unit_2_reset),
    .io_theta(cordic_unit_2_io_theta),
    .io_sin(cordic_unit_2_io_sin),
    .io_cos(cordic_unit_2_io_cos)
  );
  cordic_sin_cos_expand cordic_unit_3 ( // @[Cordic_CR.scala 271:29]
    .clock(cordic_unit_3_clock),
    .reset(cordic_unit_3_reset),
    .io_theta(cordic_unit_3_io_theta),
    .io_sin(cordic_unit_3_io_sin),
    .io_cos(cordic_unit_3_io_cos)
  );
  kronecker_v1 unit ( // @[Kronecker_V1.scala 92:22]
    .io_matrixA_1_re(unit_io_matrixA_1_re),
    .io_matrixA_1_im(unit_io_matrixA_1_im),
    .io_matrixB_1_re(unit_io_matrixB_1_re),
    .io_matrixB_1_im(unit_io_matrixB_1_im),
    .io_matrixOut_0_re(unit_io_matrixOut_0_re),
    .io_matrixOut_0_im(unit_io_matrixOut_0_im),
    .io_matrixOut_1_re(unit_io_matrixOut_1_re),
    .io_matrixOut_1_im(unit_io_matrixOut_1_im),
    .io_matrixOut_2_re(unit_io_matrixOut_2_re),
    .io_matrixOut_2_im(unit_io_matrixOut_2_im),
    .io_matrixOut_3_re(unit_io_matrixOut_3_re),
    .io_matrixOut_3_im(unit_io_matrixOut_3_im)
  );
  assign io_matrixOut_0_re = unit_io_matrixOut_0_re; // @[Space_Time_Steering_Vector.scala 88:16]
  assign io_matrixOut_0_im = unit_io_matrixOut_0_im; // @[Space_Time_Steering_Vector.scala 88:16]
  assign io_matrixOut_1_re = unit_io_matrixOut_1_re; // @[Space_Time_Steering_Vector.scala 88:16]
  assign io_matrixOut_1_im = unit_io_matrixOut_1_im; // @[Space_Time_Steering_Vector.scala 88:16]
  assign io_matrixOut_2_re = unit_io_matrixOut_2_re; // @[Space_Time_Steering_Vector.scala 88:16]
  assign io_matrixOut_2_im = unit_io_matrixOut_2_im; // @[Space_Time_Steering_Vector.scala 88:16]
  assign io_matrixOut_3_re = unit_io_matrixOut_3_re; // @[Space_Time_Steering_Vector.scala 88:16]
  assign io_matrixOut_3_im = unit_io_matrixOut_3_im; // @[Space_Time_Steering_Vector.scala 88:16]
  assign cordic_unit_clock = clock;
  assign cordic_unit_reset = reset;
  assign cordic_unit_io_theta = io_theta; // @[Cordic_CR.scala 172:26]
  assign cordic_unit_1_clock = clock;
  assign cordic_unit_1_reset = reset;
  assign cordic_unit_1_io_theta = io_psi; // @[Cordic_CR.scala 172:26]
  assign lambda_divide_divide_clock = clock;
  assign lambda_divide_divide_reset = reset;
  assign lambda_divide_divide_io_x = io_lambda; // @[Cordic_LV.scala 212:17]
  assign lambda_divide_divide_io_y = 64'sh100000000; // @[Cordic_LV.scala 213:17]
  assign cordic_unit_2_clock = clock;
  assign cordic_unit_2_reset = reset;
  assign cordic_unit_2_io_theta = _GEN_4[63:0]; // @[Cordic_CR.scala 272:26]
  assign cordic_unit_3_clock = clock;
  assign cordic_unit_3_reset = reset;
  assign cordic_unit_3_io_theta = _GEN_6[63:0]; // @[Cordic_CR.scala 272:26]
  assign unit_io_matrixA_1_re = cordic_unit_2_io_cos; // @[Space_Time_Steering_Vector.scala 65:16 76:14]
  assign unit_io_matrixA_1_im = cordic_unit_2_io_sin; // @[Space_Time_Steering_Vector.scala 65:16 77:14]
  assign unit_io_matrixB_1_re = cordic_unit_3_io_cos; // @[Space_Time_Steering_Vector.scala 66:16 83:14]
  assign unit_io_matrixB_1_im = cordic_unit_3_io_sin; // @[Space_Time_Steering_Vector.scala 66:16 84:14]
  always @(posedge clock) begin
    if (reset) begin // @[Space_Time_Steering_Vector.scala 40:39]
      reg_d_0 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 40:39]
    end else begin
      reg_d_0 <= io_d; // @[Space_Time_Steering_Vector.scala 45:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 40:39]
      reg_d_1 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 40:39]
    end else begin
      reg_d_1 <= reg_d_0; // @[Space_Time_Steering_Vector.scala 49:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 40:39]
      reg_d_2 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 40:39]
    end else begin
      reg_d_2 <= reg_d_1; // @[Space_Time_Steering_Vector.scala 49:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 40:39]
      reg_d_3 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 40:39]
    end else begin
      reg_d_3 <= reg_d_2; // @[Space_Time_Steering_Vector.scala 49:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 40:39]
      reg_d_4 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 40:39]
    end else begin
      reg_d_4 <= reg_d_3; // @[Space_Time_Steering_Vector.scala 49:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 40:39]
      reg_d_5 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 40:39]
    end else begin
      reg_d_5 <= reg_d_4; // @[Space_Time_Steering_Vector.scala 49:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 40:39]
      reg_d_6 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 40:39]
    end else begin
      reg_d_6 <= reg_d_5; // @[Space_Time_Steering_Vector.scala 49:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 40:39]
      reg_d_7 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 40:39]
    end else begin
      reg_d_7 <= reg_d_6; // @[Space_Time_Steering_Vector.scala 49:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 40:39]
      reg_d_8 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 40:39]
    end else begin
      reg_d_8 <= reg_d_7; // @[Space_Time_Steering_Vector.scala 49:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 40:39]
      reg_d_9 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 40:39]
    end else begin
      reg_d_9 <= reg_d_8; // @[Space_Time_Steering_Vector.scala 49:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 40:39]
      reg_d_10 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 40:39]
    end else begin
      reg_d_10 <= reg_d_9; // @[Space_Time_Steering_Vector.scala 49:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 40:39]
      reg_d_11 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 40:39]
    end else begin
      reg_d_11 <= reg_d_10; // @[Space_Time_Steering_Vector.scala 49:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 40:39]
      reg_d_12 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 40:39]
    end else begin
      reg_d_12 <= reg_d_11; // @[Space_Time_Steering_Vector.scala 49:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 40:39]
      reg_d_13 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 40:39]
    end else begin
      reg_d_13 <= reg_d_12; // @[Space_Time_Steering_Vector.scala 49:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 40:39]
      reg_d_14 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 40:39]
    end else begin
      reg_d_14 <= reg_d_13; // @[Space_Time_Steering_Vector.scala 49:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 41:39]
      reg_v_0 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 41:39]
    end else begin
      reg_v_0 <= io_v; // @[Space_Time_Steering_Vector.scala 46:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 41:39]
      reg_v_1 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 41:39]
    end else begin
      reg_v_1 <= reg_v_0; // @[Space_Time_Steering_Vector.scala 50:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 41:39]
      reg_v_2 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 41:39]
    end else begin
      reg_v_2 <= reg_v_1; // @[Space_Time_Steering_Vector.scala 50:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 41:39]
      reg_v_3 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 41:39]
    end else begin
      reg_v_3 <= reg_v_2; // @[Space_Time_Steering_Vector.scala 50:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 41:39]
      reg_v_4 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 41:39]
    end else begin
      reg_v_4 <= reg_v_3; // @[Space_Time_Steering_Vector.scala 50:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 41:39]
      reg_v_5 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 41:39]
    end else begin
      reg_v_5 <= reg_v_4; // @[Space_Time_Steering_Vector.scala 50:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 41:39]
      reg_v_6 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 41:39]
    end else begin
      reg_v_6 <= reg_v_5; // @[Space_Time_Steering_Vector.scala 50:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 41:39]
      reg_v_7 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 41:39]
    end else begin
      reg_v_7 <= reg_v_6; // @[Space_Time_Steering_Vector.scala 50:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 41:39]
      reg_v_8 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 41:39]
    end else begin
      reg_v_8 <= reg_v_7; // @[Space_Time_Steering_Vector.scala 50:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 41:39]
      reg_v_9 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 41:39]
    end else begin
      reg_v_9 <= reg_v_8; // @[Space_Time_Steering_Vector.scala 50:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 41:39]
      reg_v_10 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 41:39]
    end else begin
      reg_v_10 <= reg_v_9; // @[Space_Time_Steering_Vector.scala 50:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 41:39]
      reg_v_11 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 41:39]
    end else begin
      reg_v_11 <= reg_v_10; // @[Space_Time_Steering_Vector.scala 50:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 41:39]
      reg_v_12 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 41:39]
    end else begin
      reg_v_12 <= reg_v_11; // @[Space_Time_Steering_Vector.scala 50:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 41:39]
      reg_v_13 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 41:39]
    end else begin
      reg_v_13 <= reg_v_12; // @[Space_Time_Steering_Vector.scala 50:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 41:39]
      reg_v_14 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 41:39]
    end else begin
      reg_v_14 <= reg_v_13; // @[Space_Time_Steering_Vector.scala 50:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 42:39]
      reg_T_0 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 42:39]
    end else begin
      reg_T_0 <= io_T; // @[Space_Time_Steering_Vector.scala 47:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 42:39]
      reg_T_1 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 42:39]
    end else begin
      reg_T_1 <= reg_T_0; // @[Space_Time_Steering_Vector.scala 51:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 42:39]
      reg_T_2 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 42:39]
    end else begin
      reg_T_2 <= reg_T_1; // @[Space_Time_Steering_Vector.scala 51:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 42:39]
      reg_T_3 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 42:39]
    end else begin
      reg_T_3 <= reg_T_2; // @[Space_Time_Steering_Vector.scala 51:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 42:39]
      reg_T_4 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 42:39]
    end else begin
      reg_T_4 <= reg_T_3; // @[Space_Time_Steering_Vector.scala 51:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 42:39]
      reg_T_5 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 42:39]
    end else begin
      reg_T_5 <= reg_T_4; // @[Space_Time_Steering_Vector.scala 51:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 42:39]
      reg_T_6 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 42:39]
    end else begin
      reg_T_6 <= reg_T_5; // @[Space_Time_Steering_Vector.scala 51:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 42:39]
      reg_T_7 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 42:39]
    end else begin
      reg_T_7 <= reg_T_6; // @[Space_Time_Steering_Vector.scala 51:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 42:39]
      reg_T_8 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 42:39]
    end else begin
      reg_T_8 <= reg_T_7; // @[Space_Time_Steering_Vector.scala 51:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 42:39]
      reg_T_9 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 42:39]
    end else begin
      reg_T_9 <= reg_T_8; // @[Space_Time_Steering_Vector.scala 51:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 42:39]
      reg_T_10 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 42:39]
    end else begin
      reg_T_10 <= reg_T_9; // @[Space_Time_Steering_Vector.scala 51:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 42:39]
      reg_T_11 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 42:39]
    end else begin
      reg_T_11 <= reg_T_10; // @[Space_Time_Steering_Vector.scala 51:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 42:39]
      reg_T_12 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 42:39]
    end else begin
      reg_T_12 <= reg_T_11; // @[Space_Time_Steering_Vector.scala 51:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 42:39]
      reg_T_13 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 42:39]
    end else begin
      reg_T_13 <= reg_T_12; // @[Space_Time_Steering_Vector.scala 51:16]
    end
    if (reset) begin // @[Space_Time_Steering_Vector.scala 42:39]
      reg_T_14 <= 64'sh0; // @[Space_Time_Steering_Vector.scala 42:39]
    end else begin
      reg_T_14 <= reg_T_13; // @[Space_Time_Steering_Vector.scala 51:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  reg_d_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  reg_d_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  reg_d_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  reg_d_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  reg_d_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  reg_d_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  reg_d_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  reg_d_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  reg_d_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  reg_d_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  reg_d_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  reg_d_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  reg_d_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  reg_d_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  reg_d_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  reg_v_0 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  reg_v_1 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  reg_v_2 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  reg_v_3 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  reg_v_4 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  reg_v_5 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  reg_v_6 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  reg_v_7 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  reg_v_8 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  reg_v_9 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  reg_v_10 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  reg_v_11 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  reg_v_12 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  reg_v_13 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  reg_v_14 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  reg_T_0 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  reg_T_1 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  reg_T_2 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  reg_T_3 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  reg_T_4 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  reg_T_5 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  reg_T_6 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  reg_T_7 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  reg_T_8 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  reg_T_9 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  reg_T_10 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  reg_T_11 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  reg_T_12 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  reg_T_13 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  reg_T_14 = _RAND_44[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ComplexAdd(
  input  [63:0] io_op1_re,
  input  [63:0] io_op1_im,
  input  [63:0] io_op2_re,
  input  [63:0] io_op2_im,
  output [63:0] io_res_re,
  output [63:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) + $signed(io_op2_re); // @[Complex_Operater.scala 7:26]
  assign io_res_im = $signed(io_op1_im) + $signed(io_op2_im); // @[Complex_Operater.scala 8:26]
endmodule
module PE(
  input         clock,
  input         io_reset,
  input  [63:0] io_in_x_re,
  input  [63:0] io_in_x_im,
  input  [63:0] io_in_y_re,
  input  [63:0] io_in_y_im,
  output [63:0] io_out_pe_re,
  output [63:0] io_out_pe_im,
  output [63:0] io_out_x_re,
  output [63:0] io_out_x_im,
  output [63:0] io_out_y_re,
  output [63:0] io_out_y_im
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] pe_reg_mul_io_op1_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] pe_reg_mul_io_op1_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] pe_reg_mul_io_op2_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] pe_reg_mul_io_op2_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] pe_reg_mul_io_res_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] pe_reg_mul_io_res_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] pe_reg_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] pe_reg_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] pe_reg_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] pe_reg_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] pe_reg_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] pe_reg_add_io_res_im; // @[Complex_Operater.scala 13:21]
  reg [63:0] pe_reg_re; // @[Matrix_Mul_V1.scala 29:28]
  reg [63:0] pe_reg_im; // @[Matrix_Mul_V1.scala 29:28]
  reg [63:0] x_reg_re; // @[Matrix_Mul_V1.scala 30:27]
  reg [63:0] x_reg_im; // @[Matrix_Mul_V1.scala 30:27]
  reg [63:0] y_reg_re; // @[Matrix_Mul_V1.scala 31:27]
  reg [63:0] y_reg_im; // @[Matrix_Mul_V1.scala 31:27]
  ComplexMul pe_reg_mul ( // @[Complex_Operater.scala 47:21]
    .io_op1_re(pe_reg_mul_io_op1_re),
    .io_op1_im(pe_reg_mul_io_op1_im),
    .io_op2_re(pe_reg_mul_io_op2_re),
    .io_op2_im(pe_reg_mul_io_op2_im),
    .io_res_re(pe_reg_mul_io_res_re),
    .io_res_im(pe_reg_mul_io_res_im)
  );
  ComplexAdd pe_reg_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(pe_reg_add_io_op1_re),
    .io_op1_im(pe_reg_add_io_op1_im),
    .io_op2_re(pe_reg_add_io_op2_re),
    .io_op2_im(pe_reg_add_io_op2_im),
    .io_res_re(pe_reg_add_io_res_re),
    .io_res_im(pe_reg_add_io_res_im)
  );
  assign io_out_pe_re = pe_reg_re; // @[Matrix_Mul_V1.scala 50:13]
  assign io_out_pe_im = pe_reg_im; // @[Matrix_Mul_V1.scala 50:13]
  assign io_out_x_re = x_reg_re; // @[Matrix_Mul_V1.scala 51:12]
  assign io_out_x_im = x_reg_im; // @[Matrix_Mul_V1.scala 51:12]
  assign io_out_y_re = y_reg_re; // @[Matrix_Mul_V1.scala 52:12]
  assign io_out_y_im = y_reg_im; // @[Matrix_Mul_V1.scala 52:12]
  assign pe_reg_mul_io_op1_re = io_in_x_re; // @[Complex_Operater.scala 48:16]
  assign pe_reg_mul_io_op1_im = io_in_x_im; // @[Complex_Operater.scala 48:16]
  assign pe_reg_mul_io_op2_re = io_in_y_re; // @[Complex_Operater.scala 49:16]
  assign pe_reg_mul_io_op2_im = io_in_y_im; // @[Complex_Operater.scala 49:16]
  assign pe_reg_add_io_op1_re = pe_reg_re; // @[Complex_Operater.scala 14:16]
  assign pe_reg_add_io_op1_im = pe_reg_im; // @[Complex_Operater.scala 14:16]
  assign pe_reg_add_io_op2_re = pe_reg_mul_io_res_re; // @[Complex_Operater.scala 15:16]
  assign pe_reg_add_io_op2_im = pe_reg_mul_io_res_im; // @[Complex_Operater.scala 15:16]
  always @(posedge clock) begin
    if (io_reset) begin // @[Matrix_Mul_V1.scala 33:18]
      pe_reg_re <= 64'sh0; // @[Matrix_Mul_V1.scala 35:15]
    end else begin
      pe_reg_re <= pe_reg_add_io_res_re; // @[Matrix_Mul_V1.scala 43:12]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 33:18]
      pe_reg_im <= 64'sh0; // @[Matrix_Mul_V1.scala 36:15]
    end else begin
      pe_reg_im <= pe_reg_add_io_res_im; // @[Matrix_Mul_V1.scala 43:12]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 33:18]
      x_reg_re <= 64'sh0; // @[Matrix_Mul_V1.scala 37:14]
    end else begin
      x_reg_re <= io_in_x_re; // @[Matrix_Mul_V1.scala 45:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 33:18]
      x_reg_im <= 64'sh0; // @[Matrix_Mul_V1.scala 38:14]
    end else begin
      x_reg_im <= io_in_x_im; // @[Matrix_Mul_V1.scala 45:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 33:18]
      y_reg_re <= 64'sh0; // @[Matrix_Mul_V1.scala 39:14]
    end else begin
      y_reg_re <= io_in_y_re; // @[Matrix_Mul_V1.scala 46:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 33:18]
      y_reg_im <= 64'sh0; // @[Matrix_Mul_V1.scala 40:14]
    end else begin
      y_reg_im <= io_in_y_im; // @[Matrix_Mul_V1.scala 46:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pe_reg_re = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  pe_reg_im = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  x_reg_re = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  x_reg_im = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  y_reg_re = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  y_reg_im = _RAND_5[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module matrix_mul_v1(
  input         clock,
  input         io_reset,
  input         io_ready,
  input  [63:0] io_matrixA_0_re,
  input  [63:0] io_matrixA_0_im,
  input  [63:0] io_matrixA_1_re,
  input  [63:0] io_matrixA_1_im,
  input  [63:0] io_matrixA_2_re,
  input  [63:0] io_matrixA_2_im,
  input  [63:0] io_matrixA_3_re,
  input  [63:0] io_matrixA_3_im,
  input  [63:0] io_matrixB_0_re,
  input  [63:0] io_matrixB_0_im,
  input  [63:0] io_matrixB_1_re,
  input  [63:0] io_matrixB_1_im,
  input  [63:0] io_matrixB_2_re,
  input  [63:0] io_matrixB_2_im,
  input  [63:0] io_matrixB_3_re,
  input  [63:0] io_matrixB_3_im,
  output [63:0] io_matrixC_0_re,
  output [63:0] io_matrixC_0_im,
  output [63:0] io_matrixC_1_re,
  output [63:0] io_matrixC_1_im,
  output [63:0] io_matrixC_2_re,
  output [63:0] io_matrixC_2_im,
  output [63:0] io_matrixC_3_re,
  output [63:0] io_matrixC_3_im,
  output [63:0] io_matrixC_4_re,
  output [63:0] io_matrixC_4_im,
  output [63:0] io_matrixC_5_re,
  output [63:0] io_matrixC_5_im,
  output [63:0] io_matrixC_6_re,
  output [63:0] io_matrixC_6_im,
  output [63:0] io_matrixC_7_re,
  output [63:0] io_matrixC_7_im,
  output [63:0] io_matrixC_8_re,
  output [63:0] io_matrixC_8_im,
  output [63:0] io_matrixC_9_re,
  output [63:0] io_matrixC_9_im,
  output [63:0] io_matrixC_10_re,
  output [63:0] io_matrixC_10_im,
  output [63:0] io_matrixC_11_re,
  output [63:0] io_matrixC_11_im,
  output [63:0] io_matrixC_12_re,
  output [63:0] io_matrixC_12_im,
  output [63:0] io_matrixC_13_re,
  output [63:0] io_matrixC_13_im,
  output [63:0] io_matrixC_14_re,
  output [63:0] io_matrixC_14_im,
  output [63:0] io_matrixC_15_re,
  output [63:0] io_matrixC_15_im,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  PE_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_1_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_1_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_2_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_2_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_3_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_3_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_4_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_4_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_5_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_5_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_6_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_6_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_7_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_7_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_8_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_8_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_9_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_9_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_10_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_10_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_11_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_11_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_12_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_12_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_13_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_13_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_14_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_14_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_15_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_15_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  reg [63:0] regsA_0_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_0_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_1_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_1_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_2_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_2_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_3_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_3_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsB_0_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_0_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_1_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_1_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_2_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_2_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_3_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_3_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [4:0] input_point; // @[Matrix_Mul_V1.scala 84:30]
  wire [4:0] _input_point_T_1 = input_point + 5'h1; // @[Matrix_Mul_V1.scala 116:32]
  wire  _T = input_point < 5'h4; // @[Matrix_Mul_V1.scala 145:20]
  wire [3:0] _T_1 = 1'h0 * 3'h4; // @[Matrix_Mul_V1.scala 148:44]
  wire [4:0] _GEN_309 = {{1'd0}, _T_1}; // @[Matrix_Mul_V1.scala 148:60]
  wire [4:0] _T_3 = _GEN_309 + input_point; // @[Matrix_Mul_V1.scala 148:60]
  wire [63:0] _GEN_37 = 4'h1 == _T_3[3:0] ? $signed(64'sh0) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_38 = 4'h2 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_37); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_39 = 4'h3 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_38); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_40 = 4'h4 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_39); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_41 = 4'h5 == _T_3[3:0] ? $signed(regsA_1_im) : $signed(_GEN_40); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_42 = 4'h6 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_41); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_43 = 4'h7 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_42); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_44 = 4'h8 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_43); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_45 = 4'h9 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_44); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_46 = 4'ha == _T_3[3:0] ? $signed(regsA_2_im) : $signed(_GEN_45); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_47 = 4'hb == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_46); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_48 = 4'hc == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_47); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_49 = 4'hd == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_48); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_50 = 4'he == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_49); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_51 = 4'hf == _T_3[3:0] ? $signed(regsA_3_im) : $signed(_GEN_50); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_53 = 4'h1 == _T_3[3:0] ? $signed(64'sh0) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_54 = 4'h2 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_53); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_55 = 4'h3 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_54); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_56 = 4'h4 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_55); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_57 = 4'h5 == _T_3[3:0] ? $signed(regsA_1_re) : $signed(_GEN_56); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_58 = 4'h6 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_57); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_59 = 4'h7 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_58); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_60 = 4'h8 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_59); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_61 = 4'h9 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_60); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_62 = 4'ha == _T_3[3:0] ? $signed(regsA_2_re) : $signed(_GEN_61); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_63 = 4'hb == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_62); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_64 = 4'hc == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_63); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_65 = 4'hd == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_64); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_66 = 4'he == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_65); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_67 = 4'hf == _T_3[3:0] ? $signed(regsA_3_re) : $signed(_GEN_66); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [3:0] _T_5 = 1'h1 * 3'h4; // @[Matrix_Mul_V1.scala 148:44]
  wire [4:0] _GEN_310 = {{1'd0}, _T_5}; // @[Matrix_Mul_V1.scala 148:60]
  wire [4:0] _T_7 = _GEN_310 + input_point; // @[Matrix_Mul_V1.scala 148:60]
  wire [63:0] _GEN_69 = 4'h1 == _T_7[3:0] ? $signed(64'sh0) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_70 = 4'h2 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_69); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_71 = 4'h3 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_70); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_72 = 4'h4 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_71); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_73 = 4'h5 == _T_7[3:0] ? $signed(regsA_1_im) : $signed(_GEN_72); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_74 = 4'h6 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_73); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_75 = 4'h7 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_74); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_76 = 4'h8 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_75); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_77 = 4'h9 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_76); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_78 = 4'ha == _T_7[3:0] ? $signed(regsA_2_im) : $signed(_GEN_77); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_79 = 4'hb == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_78); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_80 = 4'hc == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_79); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_81 = 4'hd == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_80); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_82 = 4'he == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_81); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_83 = 4'hf == _T_7[3:0] ? $signed(regsA_3_im) : $signed(_GEN_82); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_85 = 4'h1 == _T_7[3:0] ? $signed(64'sh0) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_86 = 4'h2 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_85); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_87 = 4'h3 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_86); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_88 = 4'h4 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_87); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_89 = 4'h5 == _T_7[3:0] ? $signed(regsA_1_re) : $signed(_GEN_88); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_90 = 4'h6 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_89); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_91 = 4'h7 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_90); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_92 = 4'h8 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_91); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_93 = 4'h9 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_92); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_94 = 4'ha == _T_7[3:0] ? $signed(regsA_2_re) : $signed(_GEN_93); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_95 = 4'hb == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_94); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_96 = 4'hc == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_95); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_97 = 4'hd == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_96); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_98 = 4'he == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_97); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_99 = 4'hf == _T_7[3:0] ? $signed(regsA_3_re) : $signed(_GEN_98); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [4:0] _T_9 = 2'h2 * 3'h4; // @[Matrix_Mul_V1.scala 148:44]
  wire [4:0] _T_11 = _T_9 + input_point; // @[Matrix_Mul_V1.scala 148:60]
  wire [63:0] _GEN_101 = 4'h1 == _T_11[3:0] ? $signed(64'sh0) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_102 = 4'h2 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_101); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_103 = 4'h3 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_102); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_104 = 4'h4 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_103); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_105 = 4'h5 == _T_11[3:0] ? $signed(regsA_1_im) : $signed(_GEN_104); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_106 = 4'h6 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_105); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_107 = 4'h7 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_106); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_108 = 4'h8 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_107); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_109 = 4'h9 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_108); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_110 = 4'ha == _T_11[3:0] ? $signed(regsA_2_im) : $signed(_GEN_109); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_111 = 4'hb == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_110); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_112 = 4'hc == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_111); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_113 = 4'hd == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_112); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_114 = 4'he == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_113); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_115 = 4'hf == _T_11[3:0] ? $signed(regsA_3_im) : $signed(_GEN_114); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_117 = 4'h1 == _T_11[3:0] ? $signed(64'sh0) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_118 = 4'h2 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_117); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_119 = 4'h3 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_118); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_120 = 4'h4 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_119); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_121 = 4'h5 == _T_11[3:0] ? $signed(regsA_1_re) : $signed(_GEN_120); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_122 = 4'h6 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_121); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_123 = 4'h7 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_122); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_124 = 4'h8 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_123); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_125 = 4'h9 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_124); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_126 = 4'ha == _T_11[3:0] ? $signed(regsA_2_re) : $signed(_GEN_125); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_127 = 4'hb == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_126); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_128 = 4'hc == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_127); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_129 = 4'hd == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_128); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_130 = 4'he == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_129); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_131 = 4'hf == _T_11[3:0] ? $signed(regsA_3_re) : $signed(_GEN_130); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [4:0] _T_13 = 2'h3 * 3'h4; // @[Matrix_Mul_V1.scala 148:44]
  wire [4:0] _T_15 = _T_13 + input_point; // @[Matrix_Mul_V1.scala 148:60]
  wire [63:0] _GEN_133 = 4'h1 == _T_15[3:0] ? $signed(64'sh0) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_134 = 4'h2 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_133); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_135 = 4'h3 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_134); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_136 = 4'h4 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_135); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_137 = 4'h5 == _T_15[3:0] ? $signed(regsA_1_im) : $signed(_GEN_136); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_138 = 4'h6 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_137); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_139 = 4'h7 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_138); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_140 = 4'h8 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_139); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_141 = 4'h9 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_140); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_142 = 4'ha == _T_15[3:0] ? $signed(regsA_2_im) : $signed(_GEN_141); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_143 = 4'hb == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_142); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_144 = 4'hc == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_143); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_145 = 4'hd == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_144); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_146 = 4'he == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_145); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_147 = 4'hf == _T_15[3:0] ? $signed(regsA_3_im) : $signed(_GEN_146); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_149 = 4'h1 == _T_15[3:0] ? $signed(64'sh0) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_150 = 4'h2 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_149); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_151 = 4'h3 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_150); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_152 = 4'h4 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_151); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_153 = 4'h5 == _T_15[3:0] ? $signed(regsA_1_re) : $signed(_GEN_152); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_154 = 4'h6 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_153); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_155 = 4'h7 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_154); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_156 = 4'h8 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_155); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_157 = 4'h9 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_156); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_158 = 4'ha == _T_15[3:0] ? $signed(regsA_2_re) : $signed(_GEN_157); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_159 = 4'hb == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_158); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_160 = 4'hc == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_159); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_161 = 4'hd == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_160); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_162 = 4'he == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_161); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_163 = 4'hf == _T_15[3:0] ? $signed(regsA_3_re) : $signed(_GEN_162); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_173 = 4'h1 == _T_3[3:0] ? $signed(64'sh0) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_174 = 4'h2 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_173); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_175 = 4'h3 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_174); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_176 = 4'h4 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_175); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_177 = 4'h5 == _T_3[3:0] ? $signed(regsB_1_im) : $signed(_GEN_176); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_178 = 4'h6 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_177); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_179 = 4'h7 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_178); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_180 = 4'h8 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_179); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_181 = 4'h9 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_180); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_182 = 4'ha == _T_3[3:0] ? $signed(regsB_2_im) : $signed(_GEN_181); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_183 = 4'hb == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_182); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_184 = 4'hc == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_183); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_185 = 4'hd == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_184); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_186 = 4'he == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_185); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_187 = 4'hf == _T_3[3:0] ? $signed(regsB_3_im) : $signed(_GEN_186); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_189 = 4'h1 == _T_3[3:0] ? $signed(64'sh0) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_190 = 4'h2 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_189); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_191 = 4'h3 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_190); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_192 = 4'h4 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_191); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_193 = 4'h5 == _T_3[3:0] ? $signed(regsB_1_re) : $signed(_GEN_192); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_194 = 4'h6 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_193); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_195 = 4'h7 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_194); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_196 = 4'h8 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_195); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_197 = 4'h9 == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_196); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_198 = 4'ha == _T_3[3:0] ? $signed(regsB_2_re) : $signed(_GEN_197); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_199 = 4'hb == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_198); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_200 = 4'hc == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_199); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_201 = 4'hd == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_200); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_202 = 4'he == _T_3[3:0] ? $signed(64'sh0) : $signed(_GEN_201); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_203 = 4'hf == _T_3[3:0] ? $signed(regsB_3_re) : $signed(_GEN_202); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_205 = 4'h1 == _T_7[3:0] ? $signed(64'sh0) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_206 = 4'h2 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_205); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_207 = 4'h3 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_206); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_208 = 4'h4 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_207); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_209 = 4'h5 == _T_7[3:0] ? $signed(regsB_1_im) : $signed(_GEN_208); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_210 = 4'h6 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_209); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_211 = 4'h7 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_210); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_212 = 4'h8 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_211); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_213 = 4'h9 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_212); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_214 = 4'ha == _T_7[3:0] ? $signed(regsB_2_im) : $signed(_GEN_213); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_215 = 4'hb == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_214); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_216 = 4'hc == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_215); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_217 = 4'hd == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_216); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_218 = 4'he == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_217); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_219 = 4'hf == _T_7[3:0] ? $signed(regsB_3_im) : $signed(_GEN_218); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_221 = 4'h1 == _T_7[3:0] ? $signed(64'sh0) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_222 = 4'h2 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_221); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_223 = 4'h3 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_222); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_224 = 4'h4 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_223); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_225 = 4'h5 == _T_7[3:0] ? $signed(regsB_1_re) : $signed(_GEN_224); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_226 = 4'h6 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_225); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_227 = 4'h7 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_226); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_228 = 4'h8 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_227); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_229 = 4'h9 == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_228); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_230 = 4'ha == _T_7[3:0] ? $signed(regsB_2_re) : $signed(_GEN_229); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_231 = 4'hb == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_230); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_232 = 4'hc == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_231); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_233 = 4'hd == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_232); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_234 = 4'he == _T_7[3:0] ? $signed(64'sh0) : $signed(_GEN_233); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_235 = 4'hf == _T_7[3:0] ? $signed(regsB_3_re) : $signed(_GEN_234); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_237 = 4'h1 == _T_11[3:0] ? $signed(64'sh0) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_238 = 4'h2 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_237); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_239 = 4'h3 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_238); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_240 = 4'h4 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_239); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_241 = 4'h5 == _T_11[3:0] ? $signed(regsB_1_im) : $signed(_GEN_240); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_242 = 4'h6 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_241); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_243 = 4'h7 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_242); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_244 = 4'h8 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_243); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_245 = 4'h9 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_244); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_246 = 4'ha == _T_11[3:0] ? $signed(regsB_2_im) : $signed(_GEN_245); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_247 = 4'hb == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_246); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_248 = 4'hc == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_247); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_249 = 4'hd == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_248); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_250 = 4'he == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_249); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_251 = 4'hf == _T_11[3:0] ? $signed(regsB_3_im) : $signed(_GEN_250); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_253 = 4'h1 == _T_11[3:0] ? $signed(64'sh0) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_254 = 4'h2 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_253); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_255 = 4'h3 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_254); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_256 = 4'h4 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_255); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_257 = 4'h5 == _T_11[3:0] ? $signed(regsB_1_re) : $signed(_GEN_256); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_258 = 4'h6 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_257); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_259 = 4'h7 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_258); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_260 = 4'h8 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_259); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_261 = 4'h9 == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_260); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_262 = 4'ha == _T_11[3:0] ? $signed(regsB_2_re) : $signed(_GEN_261); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_263 = 4'hb == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_262); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_264 = 4'hc == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_263); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_265 = 4'hd == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_264); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_266 = 4'he == _T_11[3:0] ? $signed(64'sh0) : $signed(_GEN_265); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_267 = 4'hf == _T_11[3:0] ? $signed(regsB_3_re) : $signed(_GEN_266); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_269 = 4'h1 == _T_15[3:0] ? $signed(64'sh0) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_270 = 4'h2 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_269); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_271 = 4'h3 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_270); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_272 = 4'h4 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_271); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_273 = 4'h5 == _T_15[3:0] ? $signed(regsB_1_im) : $signed(_GEN_272); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_274 = 4'h6 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_273); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_275 = 4'h7 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_274); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_276 = 4'h8 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_275); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_277 = 4'h9 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_276); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_278 = 4'ha == _T_15[3:0] ? $signed(regsB_2_im) : $signed(_GEN_277); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_279 = 4'hb == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_278); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_280 = 4'hc == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_279); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_281 = 4'hd == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_280); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_282 = 4'he == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_281); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_283 = 4'hf == _T_15[3:0] ? $signed(regsB_3_im) : $signed(_GEN_282); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_285 = 4'h1 == _T_15[3:0] ? $signed(64'sh0) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_286 = 4'h2 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_285); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_287 = 4'h3 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_286); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_288 = 4'h4 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_287); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_289 = 4'h5 == _T_15[3:0] ? $signed(regsB_1_re) : $signed(_GEN_288); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_290 = 4'h6 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_289); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_291 = 4'h7 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_290); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_292 = 4'h8 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_291); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_293 = 4'h9 == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_292); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_294 = 4'ha == _T_15[3:0] ? $signed(regsB_2_re) : $signed(_GEN_293); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_295 = 4'hb == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_294); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_296 = 4'hc == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_295); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_297 = 4'hd == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_296); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_298 = 4'he == _T_15[3:0] ? $signed(64'sh0) : $signed(_GEN_297); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_299 = 4'hf == _T_15[3:0] ? $signed(regsB_3_re) : $signed(_GEN_298); // @[Matrix_Mul_V1.scala 162:{19,19}]
  PE PE ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_clock),
    .io_reset(PE_io_reset),
    .io_in_x_re(PE_io_in_x_re),
    .io_in_x_im(PE_io_in_x_im),
    .io_in_y_re(PE_io_in_y_re),
    .io_in_y_im(PE_io_in_y_im),
    .io_out_pe_re(PE_io_out_pe_re),
    .io_out_pe_im(PE_io_out_pe_im),
    .io_out_x_re(PE_io_out_x_re),
    .io_out_x_im(PE_io_out_x_im),
    .io_out_y_re(PE_io_out_y_re),
    .io_out_y_im(PE_io_out_y_im)
  );
  PE PE_1 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_1_clock),
    .io_reset(PE_1_io_reset),
    .io_in_x_re(PE_1_io_in_x_re),
    .io_in_x_im(PE_1_io_in_x_im),
    .io_in_y_re(PE_1_io_in_y_re),
    .io_in_y_im(PE_1_io_in_y_im),
    .io_out_pe_re(PE_1_io_out_pe_re),
    .io_out_pe_im(PE_1_io_out_pe_im),
    .io_out_x_re(PE_1_io_out_x_re),
    .io_out_x_im(PE_1_io_out_x_im),
    .io_out_y_re(PE_1_io_out_y_re),
    .io_out_y_im(PE_1_io_out_y_im)
  );
  PE PE_2 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_2_clock),
    .io_reset(PE_2_io_reset),
    .io_in_x_re(PE_2_io_in_x_re),
    .io_in_x_im(PE_2_io_in_x_im),
    .io_in_y_re(PE_2_io_in_y_re),
    .io_in_y_im(PE_2_io_in_y_im),
    .io_out_pe_re(PE_2_io_out_pe_re),
    .io_out_pe_im(PE_2_io_out_pe_im),
    .io_out_x_re(PE_2_io_out_x_re),
    .io_out_x_im(PE_2_io_out_x_im),
    .io_out_y_re(PE_2_io_out_y_re),
    .io_out_y_im(PE_2_io_out_y_im)
  );
  PE PE_3 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_3_clock),
    .io_reset(PE_3_io_reset),
    .io_in_x_re(PE_3_io_in_x_re),
    .io_in_x_im(PE_3_io_in_x_im),
    .io_in_y_re(PE_3_io_in_y_re),
    .io_in_y_im(PE_3_io_in_y_im),
    .io_out_pe_re(PE_3_io_out_pe_re),
    .io_out_pe_im(PE_3_io_out_pe_im),
    .io_out_x_re(PE_3_io_out_x_re),
    .io_out_x_im(PE_3_io_out_x_im),
    .io_out_y_re(PE_3_io_out_y_re),
    .io_out_y_im(PE_3_io_out_y_im)
  );
  PE PE_4 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_4_clock),
    .io_reset(PE_4_io_reset),
    .io_in_x_re(PE_4_io_in_x_re),
    .io_in_x_im(PE_4_io_in_x_im),
    .io_in_y_re(PE_4_io_in_y_re),
    .io_in_y_im(PE_4_io_in_y_im),
    .io_out_pe_re(PE_4_io_out_pe_re),
    .io_out_pe_im(PE_4_io_out_pe_im),
    .io_out_x_re(PE_4_io_out_x_re),
    .io_out_x_im(PE_4_io_out_x_im),
    .io_out_y_re(PE_4_io_out_y_re),
    .io_out_y_im(PE_4_io_out_y_im)
  );
  PE PE_5 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_5_clock),
    .io_reset(PE_5_io_reset),
    .io_in_x_re(PE_5_io_in_x_re),
    .io_in_x_im(PE_5_io_in_x_im),
    .io_in_y_re(PE_5_io_in_y_re),
    .io_in_y_im(PE_5_io_in_y_im),
    .io_out_pe_re(PE_5_io_out_pe_re),
    .io_out_pe_im(PE_5_io_out_pe_im),
    .io_out_x_re(PE_5_io_out_x_re),
    .io_out_x_im(PE_5_io_out_x_im),
    .io_out_y_re(PE_5_io_out_y_re),
    .io_out_y_im(PE_5_io_out_y_im)
  );
  PE PE_6 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_6_clock),
    .io_reset(PE_6_io_reset),
    .io_in_x_re(PE_6_io_in_x_re),
    .io_in_x_im(PE_6_io_in_x_im),
    .io_in_y_re(PE_6_io_in_y_re),
    .io_in_y_im(PE_6_io_in_y_im),
    .io_out_pe_re(PE_6_io_out_pe_re),
    .io_out_pe_im(PE_6_io_out_pe_im),
    .io_out_x_re(PE_6_io_out_x_re),
    .io_out_x_im(PE_6_io_out_x_im),
    .io_out_y_re(PE_6_io_out_y_re),
    .io_out_y_im(PE_6_io_out_y_im)
  );
  PE PE_7 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_7_clock),
    .io_reset(PE_7_io_reset),
    .io_in_x_re(PE_7_io_in_x_re),
    .io_in_x_im(PE_7_io_in_x_im),
    .io_in_y_re(PE_7_io_in_y_re),
    .io_in_y_im(PE_7_io_in_y_im),
    .io_out_pe_re(PE_7_io_out_pe_re),
    .io_out_pe_im(PE_7_io_out_pe_im),
    .io_out_x_re(PE_7_io_out_x_re),
    .io_out_x_im(PE_7_io_out_x_im),
    .io_out_y_re(PE_7_io_out_y_re),
    .io_out_y_im(PE_7_io_out_y_im)
  );
  PE PE_8 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_8_clock),
    .io_reset(PE_8_io_reset),
    .io_in_x_re(PE_8_io_in_x_re),
    .io_in_x_im(PE_8_io_in_x_im),
    .io_in_y_re(PE_8_io_in_y_re),
    .io_in_y_im(PE_8_io_in_y_im),
    .io_out_pe_re(PE_8_io_out_pe_re),
    .io_out_pe_im(PE_8_io_out_pe_im),
    .io_out_x_re(PE_8_io_out_x_re),
    .io_out_x_im(PE_8_io_out_x_im),
    .io_out_y_re(PE_8_io_out_y_re),
    .io_out_y_im(PE_8_io_out_y_im)
  );
  PE PE_9 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_9_clock),
    .io_reset(PE_9_io_reset),
    .io_in_x_re(PE_9_io_in_x_re),
    .io_in_x_im(PE_9_io_in_x_im),
    .io_in_y_re(PE_9_io_in_y_re),
    .io_in_y_im(PE_9_io_in_y_im),
    .io_out_pe_re(PE_9_io_out_pe_re),
    .io_out_pe_im(PE_9_io_out_pe_im),
    .io_out_x_re(PE_9_io_out_x_re),
    .io_out_x_im(PE_9_io_out_x_im),
    .io_out_y_re(PE_9_io_out_y_re),
    .io_out_y_im(PE_9_io_out_y_im)
  );
  PE PE_10 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_10_clock),
    .io_reset(PE_10_io_reset),
    .io_in_x_re(PE_10_io_in_x_re),
    .io_in_x_im(PE_10_io_in_x_im),
    .io_in_y_re(PE_10_io_in_y_re),
    .io_in_y_im(PE_10_io_in_y_im),
    .io_out_pe_re(PE_10_io_out_pe_re),
    .io_out_pe_im(PE_10_io_out_pe_im),
    .io_out_x_re(PE_10_io_out_x_re),
    .io_out_x_im(PE_10_io_out_x_im),
    .io_out_y_re(PE_10_io_out_y_re),
    .io_out_y_im(PE_10_io_out_y_im)
  );
  PE PE_11 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_11_clock),
    .io_reset(PE_11_io_reset),
    .io_in_x_re(PE_11_io_in_x_re),
    .io_in_x_im(PE_11_io_in_x_im),
    .io_in_y_re(PE_11_io_in_y_re),
    .io_in_y_im(PE_11_io_in_y_im),
    .io_out_pe_re(PE_11_io_out_pe_re),
    .io_out_pe_im(PE_11_io_out_pe_im),
    .io_out_x_re(PE_11_io_out_x_re),
    .io_out_x_im(PE_11_io_out_x_im),
    .io_out_y_re(PE_11_io_out_y_re),
    .io_out_y_im(PE_11_io_out_y_im)
  );
  PE PE_12 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_12_clock),
    .io_reset(PE_12_io_reset),
    .io_in_x_re(PE_12_io_in_x_re),
    .io_in_x_im(PE_12_io_in_x_im),
    .io_in_y_re(PE_12_io_in_y_re),
    .io_in_y_im(PE_12_io_in_y_im),
    .io_out_pe_re(PE_12_io_out_pe_re),
    .io_out_pe_im(PE_12_io_out_pe_im),
    .io_out_x_re(PE_12_io_out_x_re),
    .io_out_x_im(PE_12_io_out_x_im),
    .io_out_y_re(PE_12_io_out_y_re),
    .io_out_y_im(PE_12_io_out_y_im)
  );
  PE PE_13 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_13_clock),
    .io_reset(PE_13_io_reset),
    .io_in_x_re(PE_13_io_in_x_re),
    .io_in_x_im(PE_13_io_in_x_im),
    .io_in_y_re(PE_13_io_in_y_re),
    .io_in_y_im(PE_13_io_in_y_im),
    .io_out_pe_re(PE_13_io_out_pe_re),
    .io_out_pe_im(PE_13_io_out_pe_im),
    .io_out_x_re(PE_13_io_out_x_re),
    .io_out_x_im(PE_13_io_out_x_im),
    .io_out_y_re(PE_13_io_out_y_re),
    .io_out_y_im(PE_13_io_out_y_im)
  );
  PE PE_14 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_14_clock),
    .io_reset(PE_14_io_reset),
    .io_in_x_re(PE_14_io_in_x_re),
    .io_in_x_im(PE_14_io_in_x_im),
    .io_in_y_re(PE_14_io_in_y_re),
    .io_in_y_im(PE_14_io_in_y_im),
    .io_out_pe_re(PE_14_io_out_pe_re),
    .io_out_pe_im(PE_14_io_out_pe_im),
    .io_out_x_re(PE_14_io_out_x_re),
    .io_out_x_im(PE_14_io_out_x_im),
    .io_out_y_re(PE_14_io_out_y_re),
    .io_out_y_im(PE_14_io_out_y_im)
  );
  PE PE_15 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_15_clock),
    .io_reset(PE_15_io_reset),
    .io_in_x_re(PE_15_io_in_x_re),
    .io_in_x_im(PE_15_io_in_x_im),
    .io_in_y_re(PE_15_io_in_y_re),
    .io_in_y_im(PE_15_io_in_y_im),
    .io_out_pe_re(PE_15_io_out_pe_re),
    .io_out_pe_im(PE_15_io_out_pe_im),
    .io_out_x_re(PE_15_io_out_x_re),
    .io_out_x_im(PE_15_io_out_x_im),
    .io_out_y_re(PE_15_io_out_y_re),
    .io_out_y_im(PE_15_io_out_y_im)
  );
  assign io_matrixC_0_re = PE_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_0_im = PE_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_1_re = PE_1_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_1_im = PE_1_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_2_re = PE_2_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_2_im = PE_2_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_3_re = PE_3_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_3_im = PE_3_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_4_re = PE_4_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_4_im = PE_4_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_5_re = PE_5_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_5_im = PE_5_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_6_re = PE_6_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_6_im = PE_6_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_7_re = PE_7_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_7_im = PE_7_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_8_re = PE_8_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_8_im = PE_8_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_9_re = PE_9_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_9_im = PE_9_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_10_re = PE_10_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_10_im = PE_10_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_11_re = PE_11_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_11_im = PE_11_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_12_re = PE_12_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_12_im = PE_12_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_13_re = PE_13_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_13_im = PE_13_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_14_re = PE_14_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_14_im = PE_14_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_15_re = PE_15_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_15_im = PE_15_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_valid = input_point >= 5'h7; // @[Matrix_Mul_V1.scala 188:20]
  assign PE_clock = clock;
  assign PE_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_io_in_x_re = input_point < 5'h4 ? $signed(_GEN_67) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_io_in_x_im = input_point < 5'h4 ? $signed(_GEN_51) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_io_in_y_re = _T ? $signed(_GEN_203) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_io_in_y_im = _T ? $signed(_GEN_187) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_1_clock = clock;
  assign PE_1_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_1_io_in_x_re = PE_io_out_x_re; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_1_io_in_x_im = PE_io_out_x_im; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_1_io_in_y_re = _T ? $signed(_GEN_235) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_1_io_in_y_im = _T ? $signed(_GEN_219) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_2_clock = clock;
  assign PE_2_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_2_io_in_x_re = PE_1_io_out_x_re; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_2_io_in_x_im = PE_1_io_out_x_im; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_2_io_in_y_re = _T ? $signed(_GEN_267) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_2_io_in_y_im = _T ? $signed(_GEN_251) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_3_clock = clock;
  assign PE_3_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_3_io_in_x_re = PE_2_io_out_x_re; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_3_io_in_x_im = PE_2_io_out_x_im; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_3_io_in_y_re = _T ? $signed(_GEN_299) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_3_io_in_y_im = _T ? $signed(_GEN_283) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_4_clock = clock;
  assign PE_4_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_4_io_in_x_re = input_point < 5'h4 ? $signed(_GEN_99) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_4_io_in_x_im = input_point < 5'h4 ? $signed(_GEN_83) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_4_io_in_y_re = PE_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_4_io_in_y_im = PE_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_5_clock = clock;
  assign PE_5_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_5_io_in_x_re = PE_4_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_5_io_in_x_im = PE_4_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_5_io_in_y_re = PE_1_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_5_io_in_y_im = PE_1_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_6_clock = clock;
  assign PE_6_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_6_io_in_x_re = PE_5_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_6_io_in_x_im = PE_5_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_6_io_in_y_re = PE_2_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_6_io_in_y_im = PE_2_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_7_clock = clock;
  assign PE_7_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_7_io_in_x_re = PE_6_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_7_io_in_x_im = PE_6_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_7_io_in_y_re = PE_3_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_7_io_in_y_im = PE_3_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_8_clock = clock;
  assign PE_8_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_8_io_in_x_re = input_point < 5'h4 ? $signed(_GEN_131) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_8_io_in_x_im = input_point < 5'h4 ? $signed(_GEN_115) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_8_io_in_y_re = PE_4_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_8_io_in_y_im = PE_4_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_9_clock = clock;
  assign PE_9_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_9_io_in_x_re = PE_8_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_9_io_in_x_im = PE_8_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_9_io_in_y_re = PE_5_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_9_io_in_y_im = PE_5_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_10_clock = clock;
  assign PE_10_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_10_io_in_x_re = PE_9_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_10_io_in_x_im = PE_9_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_10_io_in_y_re = PE_6_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_10_io_in_y_im = PE_6_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_11_clock = clock;
  assign PE_11_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_11_io_in_x_re = PE_10_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_11_io_in_x_im = PE_10_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_11_io_in_y_re = PE_7_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_11_io_in_y_im = PE_7_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_12_clock = clock;
  assign PE_12_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_12_io_in_x_re = input_point < 5'h4 ? $signed(_GEN_163) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_12_io_in_x_im = input_point < 5'h4 ? $signed(_GEN_147) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_12_io_in_y_re = PE_8_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_12_io_in_y_im = PE_8_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_13_clock = clock;
  assign PE_13_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_13_io_in_x_re = PE_12_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_13_io_in_x_im = PE_12_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_13_io_in_y_re = PE_9_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_13_io_in_y_im = PE_9_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_14_clock = clock;
  assign PE_14_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_14_io_in_x_re = PE_13_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_14_io_in_x_im = PE_13_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_14_io_in_y_re = PE_10_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_14_io_in_y_im = PE_10_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_15_clock = clock;
  assign PE_15_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_15_io_in_x_re = PE_14_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_15_io_in_x_im = PE_14_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_15_io_in_y_re = PE_11_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_15_io_in_y_im = PE_11_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  always @(posedge clock) begin
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_0_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_0_re <= io_matrixA_0_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_0_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_0_im <= io_matrixA_0_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_1_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_1_re <= io_matrixA_1_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_1_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_1_im <= io_matrixA_1_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_2_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_2_re <= io_matrixA_2_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_2_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_2_im <= io_matrixA_2_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_3_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_3_re <= io_matrixA_3_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_3_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_3_im <= io_matrixA_3_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_0_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_0_re <= io_matrixB_0_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_0_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_0_im <= io_matrixB_0_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_1_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_1_re <= io_matrixB_1_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_1_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_1_im <= io_matrixB_1_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_2_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_2_re <= io_matrixB_2_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_2_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_2_im <= io_matrixB_2_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_3_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_3_re <= io_matrixB_3_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_3_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_3_im <= io_matrixB_3_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      input_point <= 5'h0; // @[Matrix_Mul_V1.scala 99:17]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      input_point <= 5'h0; // @[Matrix_Mul_V1.scala 108:17]
    end else begin
      input_point <= _input_point_T_1; // @[Matrix_Mul_V1.scala 116:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regsA_0_re = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regsA_0_im = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  regsA_1_re = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  regsA_1_im = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  regsA_2_re = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  regsA_2_im = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  regsA_3_re = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  regsA_3_im = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  regsB_0_re = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  regsB_0_im = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  regsB_1_re = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  regsB_1_im = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  regsB_2_re = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  regsB_2_im = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  regsB_3_re = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  regsB_3_im = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  input_point = _RAND_16[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module complex_vector_divide_fixedPoint(
  input         clock,
  input         reset,
  input  [63:0] io_dividedVector_0_re,
  input  [63:0] io_dividedVector_0_im,
  input  [63:0] io_dividedVector_1_re,
  input  [63:0] io_dividedVector_1_im,
  input  [63:0] io_dividedVector_2_re,
  input  [63:0] io_dividedVector_2_im,
  input  [63:0] io_dividedVector_3_re,
  input  [63:0] io_dividedVector_3_im,
  input  [63:0] io_dividedVector_4_re,
  input  [63:0] io_dividedVector_4_im,
  input  [63:0] io_dividedVector_5_re,
  input  [63:0] io_dividedVector_5_im,
  input  [63:0] io_dividedVector_6_re,
  input  [63:0] io_dividedVector_6_im,
  input  [63:0] io_dividedVector_7_re,
  input  [63:0] io_dividedVector_7_im,
  input  [63:0] io_dividedVector_8_re,
  input  [63:0] io_dividedVector_8_im,
  input  [63:0] io_dividedVector_9_re,
  input  [63:0] io_dividedVector_9_im,
  input  [63:0] io_dividedVector_10_re,
  input  [63:0] io_dividedVector_10_im,
  input  [63:0] io_dividedVector_11_re,
  input  [63:0] io_dividedVector_11_im,
  input  [63:0] io_dividedVector_12_re,
  input  [63:0] io_dividedVector_12_im,
  input  [63:0] io_dividedVector_13_re,
  input  [63:0] io_dividedVector_13_im,
  input  [63:0] io_dividedVector_14_re,
  input  [63:0] io_dividedVector_14_im,
  input  [63:0] io_dividedVector_15_re,
  input  [63:0] io_dividedVector_15_im,
  output [63:0] io_vectorOut_0_re,
  output [63:0] io_vectorOut_0_im,
  output [63:0] io_vectorOut_1_re,
  output [63:0] io_vectorOut_1_im,
  output [63:0] io_vectorOut_2_re,
  output [63:0] io_vectorOut_2_im,
  output [63:0] io_vectorOut_3_re,
  output [63:0] io_vectorOut_3_im,
  output [63:0] io_vectorOut_4_re,
  output [63:0] io_vectorOut_4_im,
  output [63:0] io_vectorOut_5_re,
  output [63:0] io_vectorOut_5_im,
  output [63:0] io_vectorOut_6_re,
  output [63:0] io_vectorOut_6_im,
  output [63:0] io_vectorOut_7_re,
  output [63:0] io_vectorOut_7_im,
  output [63:0] io_vectorOut_8_re,
  output [63:0] io_vectorOut_8_im,
  output [63:0] io_vectorOut_9_re,
  output [63:0] io_vectorOut_9_im,
  output [63:0] io_vectorOut_10_re,
  output [63:0] io_vectorOut_10_im,
  output [63:0] io_vectorOut_11_re,
  output [63:0] io_vectorOut_11_im,
  output [63:0] io_vectorOut_12_re,
  output [63:0] io_vectorOut_12_im,
  output [63:0] io_vectorOut_13_re,
  output [63:0] io_vectorOut_13_im,
  output [63:0] io_vectorOut_14_re,
  output [63:0] io_vectorOut_14_im,
  output [63:0] io_vectorOut_15_re,
  output [63:0] io_vectorOut_15_im
);
  wire  io_vectorOut_0_re_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_0_re_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_0_re_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_0_re_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_0_re_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_0_im_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_0_im_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_0_im_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_0_im_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_0_im_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_1_re_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_1_re_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_1_re_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_1_re_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_1_re_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_1_im_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_1_im_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_1_im_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_1_im_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_1_im_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_2_re_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_2_re_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_2_re_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_2_re_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_2_re_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_2_im_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_2_im_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_2_im_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_2_im_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_2_im_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_3_re_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_3_re_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_3_re_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_3_re_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_3_re_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_3_im_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_3_im_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_3_im_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_3_im_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_3_im_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_4_re_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_4_re_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_4_re_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_4_re_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_4_re_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_4_im_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_4_im_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_4_im_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_4_im_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_4_im_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_5_re_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_5_re_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_5_re_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_5_re_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_5_re_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_5_im_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_5_im_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_5_im_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_5_im_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_5_im_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_6_re_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_6_re_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_6_re_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_6_re_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_6_re_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_6_im_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_6_im_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_6_im_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_6_im_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_6_im_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_7_re_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_7_re_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_7_re_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_7_re_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_7_re_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_7_im_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_7_im_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_7_im_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_7_im_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_7_im_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_8_re_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_8_re_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_8_re_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_8_re_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_8_re_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_8_im_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_8_im_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_8_im_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_8_im_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_8_im_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_9_re_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_9_re_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_9_re_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_9_re_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_9_re_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_9_im_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_9_im_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_9_im_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_9_im_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_9_im_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_10_re_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_10_re_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_10_re_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_10_re_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_10_re_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_10_im_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_10_im_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_10_im_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_10_im_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_10_im_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_11_re_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_11_re_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_11_re_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_11_re_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_11_re_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_11_im_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_11_im_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_11_im_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_11_im_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_11_im_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_12_re_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_12_re_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_12_re_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_12_re_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_12_re_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_12_im_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_12_im_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_12_im_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_12_im_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_12_im_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_13_re_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_13_re_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_13_re_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_13_re_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_13_re_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_13_im_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_13_im_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_13_im_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_13_im_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_13_im_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_14_re_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_14_re_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_14_re_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_14_re_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_14_re_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_14_im_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_14_im_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_14_im_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_14_im_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_14_im_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_15_re_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_15_re_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_15_re_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_15_re_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_15_re_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_15_im_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  io_vectorOut_15_im_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_15_im_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_15_im_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] io_vectorOut_15_im_divide_io_z; // @[Cordic_LV.scala 211:24]
  cordic_divide io_vectorOut_0_re_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_0_re_divide_clock),
    .reset(io_vectorOut_0_re_divide_reset),
    .io_x(io_vectorOut_0_re_divide_io_x),
    .io_y(io_vectorOut_0_re_divide_io_y),
    .io_z(io_vectorOut_0_re_divide_io_z)
  );
  cordic_divide io_vectorOut_0_im_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_0_im_divide_clock),
    .reset(io_vectorOut_0_im_divide_reset),
    .io_x(io_vectorOut_0_im_divide_io_x),
    .io_y(io_vectorOut_0_im_divide_io_y),
    .io_z(io_vectorOut_0_im_divide_io_z)
  );
  cordic_divide io_vectorOut_1_re_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_1_re_divide_clock),
    .reset(io_vectorOut_1_re_divide_reset),
    .io_x(io_vectorOut_1_re_divide_io_x),
    .io_y(io_vectorOut_1_re_divide_io_y),
    .io_z(io_vectorOut_1_re_divide_io_z)
  );
  cordic_divide io_vectorOut_1_im_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_1_im_divide_clock),
    .reset(io_vectorOut_1_im_divide_reset),
    .io_x(io_vectorOut_1_im_divide_io_x),
    .io_y(io_vectorOut_1_im_divide_io_y),
    .io_z(io_vectorOut_1_im_divide_io_z)
  );
  cordic_divide io_vectorOut_2_re_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_2_re_divide_clock),
    .reset(io_vectorOut_2_re_divide_reset),
    .io_x(io_vectorOut_2_re_divide_io_x),
    .io_y(io_vectorOut_2_re_divide_io_y),
    .io_z(io_vectorOut_2_re_divide_io_z)
  );
  cordic_divide io_vectorOut_2_im_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_2_im_divide_clock),
    .reset(io_vectorOut_2_im_divide_reset),
    .io_x(io_vectorOut_2_im_divide_io_x),
    .io_y(io_vectorOut_2_im_divide_io_y),
    .io_z(io_vectorOut_2_im_divide_io_z)
  );
  cordic_divide io_vectorOut_3_re_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_3_re_divide_clock),
    .reset(io_vectorOut_3_re_divide_reset),
    .io_x(io_vectorOut_3_re_divide_io_x),
    .io_y(io_vectorOut_3_re_divide_io_y),
    .io_z(io_vectorOut_3_re_divide_io_z)
  );
  cordic_divide io_vectorOut_3_im_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_3_im_divide_clock),
    .reset(io_vectorOut_3_im_divide_reset),
    .io_x(io_vectorOut_3_im_divide_io_x),
    .io_y(io_vectorOut_3_im_divide_io_y),
    .io_z(io_vectorOut_3_im_divide_io_z)
  );
  cordic_divide io_vectorOut_4_re_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_4_re_divide_clock),
    .reset(io_vectorOut_4_re_divide_reset),
    .io_x(io_vectorOut_4_re_divide_io_x),
    .io_y(io_vectorOut_4_re_divide_io_y),
    .io_z(io_vectorOut_4_re_divide_io_z)
  );
  cordic_divide io_vectorOut_4_im_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_4_im_divide_clock),
    .reset(io_vectorOut_4_im_divide_reset),
    .io_x(io_vectorOut_4_im_divide_io_x),
    .io_y(io_vectorOut_4_im_divide_io_y),
    .io_z(io_vectorOut_4_im_divide_io_z)
  );
  cordic_divide io_vectorOut_5_re_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_5_re_divide_clock),
    .reset(io_vectorOut_5_re_divide_reset),
    .io_x(io_vectorOut_5_re_divide_io_x),
    .io_y(io_vectorOut_5_re_divide_io_y),
    .io_z(io_vectorOut_5_re_divide_io_z)
  );
  cordic_divide io_vectorOut_5_im_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_5_im_divide_clock),
    .reset(io_vectorOut_5_im_divide_reset),
    .io_x(io_vectorOut_5_im_divide_io_x),
    .io_y(io_vectorOut_5_im_divide_io_y),
    .io_z(io_vectorOut_5_im_divide_io_z)
  );
  cordic_divide io_vectorOut_6_re_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_6_re_divide_clock),
    .reset(io_vectorOut_6_re_divide_reset),
    .io_x(io_vectorOut_6_re_divide_io_x),
    .io_y(io_vectorOut_6_re_divide_io_y),
    .io_z(io_vectorOut_6_re_divide_io_z)
  );
  cordic_divide io_vectorOut_6_im_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_6_im_divide_clock),
    .reset(io_vectorOut_6_im_divide_reset),
    .io_x(io_vectorOut_6_im_divide_io_x),
    .io_y(io_vectorOut_6_im_divide_io_y),
    .io_z(io_vectorOut_6_im_divide_io_z)
  );
  cordic_divide io_vectorOut_7_re_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_7_re_divide_clock),
    .reset(io_vectorOut_7_re_divide_reset),
    .io_x(io_vectorOut_7_re_divide_io_x),
    .io_y(io_vectorOut_7_re_divide_io_y),
    .io_z(io_vectorOut_7_re_divide_io_z)
  );
  cordic_divide io_vectorOut_7_im_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_7_im_divide_clock),
    .reset(io_vectorOut_7_im_divide_reset),
    .io_x(io_vectorOut_7_im_divide_io_x),
    .io_y(io_vectorOut_7_im_divide_io_y),
    .io_z(io_vectorOut_7_im_divide_io_z)
  );
  cordic_divide io_vectorOut_8_re_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_8_re_divide_clock),
    .reset(io_vectorOut_8_re_divide_reset),
    .io_x(io_vectorOut_8_re_divide_io_x),
    .io_y(io_vectorOut_8_re_divide_io_y),
    .io_z(io_vectorOut_8_re_divide_io_z)
  );
  cordic_divide io_vectorOut_8_im_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_8_im_divide_clock),
    .reset(io_vectorOut_8_im_divide_reset),
    .io_x(io_vectorOut_8_im_divide_io_x),
    .io_y(io_vectorOut_8_im_divide_io_y),
    .io_z(io_vectorOut_8_im_divide_io_z)
  );
  cordic_divide io_vectorOut_9_re_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_9_re_divide_clock),
    .reset(io_vectorOut_9_re_divide_reset),
    .io_x(io_vectorOut_9_re_divide_io_x),
    .io_y(io_vectorOut_9_re_divide_io_y),
    .io_z(io_vectorOut_9_re_divide_io_z)
  );
  cordic_divide io_vectorOut_9_im_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_9_im_divide_clock),
    .reset(io_vectorOut_9_im_divide_reset),
    .io_x(io_vectorOut_9_im_divide_io_x),
    .io_y(io_vectorOut_9_im_divide_io_y),
    .io_z(io_vectorOut_9_im_divide_io_z)
  );
  cordic_divide io_vectorOut_10_re_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_10_re_divide_clock),
    .reset(io_vectorOut_10_re_divide_reset),
    .io_x(io_vectorOut_10_re_divide_io_x),
    .io_y(io_vectorOut_10_re_divide_io_y),
    .io_z(io_vectorOut_10_re_divide_io_z)
  );
  cordic_divide io_vectorOut_10_im_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_10_im_divide_clock),
    .reset(io_vectorOut_10_im_divide_reset),
    .io_x(io_vectorOut_10_im_divide_io_x),
    .io_y(io_vectorOut_10_im_divide_io_y),
    .io_z(io_vectorOut_10_im_divide_io_z)
  );
  cordic_divide io_vectorOut_11_re_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_11_re_divide_clock),
    .reset(io_vectorOut_11_re_divide_reset),
    .io_x(io_vectorOut_11_re_divide_io_x),
    .io_y(io_vectorOut_11_re_divide_io_y),
    .io_z(io_vectorOut_11_re_divide_io_z)
  );
  cordic_divide io_vectorOut_11_im_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_11_im_divide_clock),
    .reset(io_vectorOut_11_im_divide_reset),
    .io_x(io_vectorOut_11_im_divide_io_x),
    .io_y(io_vectorOut_11_im_divide_io_y),
    .io_z(io_vectorOut_11_im_divide_io_z)
  );
  cordic_divide io_vectorOut_12_re_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_12_re_divide_clock),
    .reset(io_vectorOut_12_re_divide_reset),
    .io_x(io_vectorOut_12_re_divide_io_x),
    .io_y(io_vectorOut_12_re_divide_io_y),
    .io_z(io_vectorOut_12_re_divide_io_z)
  );
  cordic_divide io_vectorOut_12_im_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_12_im_divide_clock),
    .reset(io_vectorOut_12_im_divide_reset),
    .io_x(io_vectorOut_12_im_divide_io_x),
    .io_y(io_vectorOut_12_im_divide_io_y),
    .io_z(io_vectorOut_12_im_divide_io_z)
  );
  cordic_divide io_vectorOut_13_re_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_13_re_divide_clock),
    .reset(io_vectorOut_13_re_divide_reset),
    .io_x(io_vectorOut_13_re_divide_io_x),
    .io_y(io_vectorOut_13_re_divide_io_y),
    .io_z(io_vectorOut_13_re_divide_io_z)
  );
  cordic_divide io_vectorOut_13_im_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_13_im_divide_clock),
    .reset(io_vectorOut_13_im_divide_reset),
    .io_x(io_vectorOut_13_im_divide_io_x),
    .io_y(io_vectorOut_13_im_divide_io_y),
    .io_z(io_vectorOut_13_im_divide_io_z)
  );
  cordic_divide io_vectorOut_14_re_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_14_re_divide_clock),
    .reset(io_vectorOut_14_re_divide_reset),
    .io_x(io_vectorOut_14_re_divide_io_x),
    .io_y(io_vectorOut_14_re_divide_io_y),
    .io_z(io_vectorOut_14_re_divide_io_z)
  );
  cordic_divide io_vectorOut_14_im_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_14_im_divide_clock),
    .reset(io_vectorOut_14_im_divide_reset),
    .io_x(io_vectorOut_14_im_divide_io_x),
    .io_y(io_vectorOut_14_im_divide_io_y),
    .io_z(io_vectorOut_14_im_divide_io_z)
  );
  cordic_divide io_vectorOut_15_re_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_15_re_divide_clock),
    .reset(io_vectorOut_15_re_divide_reset),
    .io_x(io_vectorOut_15_re_divide_io_x),
    .io_y(io_vectorOut_15_re_divide_io_y),
    .io_z(io_vectorOut_15_re_divide_io_z)
  );
  cordic_divide io_vectorOut_15_im_divide ( // @[Cordic_LV.scala 211:24]
    .clock(io_vectorOut_15_im_divide_clock),
    .reset(io_vectorOut_15_im_divide_reset),
    .io_x(io_vectorOut_15_im_divide_io_x),
    .io_y(io_vectorOut_15_im_divide_io_y),
    .io_z(io_vectorOut_15_im_divide_io_z)
  );
  assign io_vectorOut_0_re = io_vectorOut_0_re_divide_io_z; // @[Complex_Vector_Divide.scala 43:24]
  assign io_vectorOut_0_im = io_vectorOut_0_im_divide_io_z; // @[Complex_Vector_Divide.scala 44:24]
  assign io_vectorOut_1_re = io_vectorOut_1_re_divide_io_z; // @[Complex_Vector_Divide.scala 43:24]
  assign io_vectorOut_1_im = io_vectorOut_1_im_divide_io_z; // @[Complex_Vector_Divide.scala 44:24]
  assign io_vectorOut_2_re = io_vectorOut_2_re_divide_io_z; // @[Complex_Vector_Divide.scala 43:24]
  assign io_vectorOut_2_im = io_vectorOut_2_im_divide_io_z; // @[Complex_Vector_Divide.scala 44:24]
  assign io_vectorOut_3_re = io_vectorOut_3_re_divide_io_z; // @[Complex_Vector_Divide.scala 43:24]
  assign io_vectorOut_3_im = io_vectorOut_3_im_divide_io_z; // @[Complex_Vector_Divide.scala 44:24]
  assign io_vectorOut_4_re = io_vectorOut_4_re_divide_io_z; // @[Complex_Vector_Divide.scala 43:24]
  assign io_vectorOut_4_im = io_vectorOut_4_im_divide_io_z; // @[Complex_Vector_Divide.scala 44:24]
  assign io_vectorOut_5_re = io_vectorOut_5_re_divide_io_z; // @[Complex_Vector_Divide.scala 43:24]
  assign io_vectorOut_5_im = io_vectorOut_5_im_divide_io_z; // @[Complex_Vector_Divide.scala 44:24]
  assign io_vectorOut_6_re = io_vectorOut_6_re_divide_io_z; // @[Complex_Vector_Divide.scala 43:24]
  assign io_vectorOut_6_im = io_vectorOut_6_im_divide_io_z; // @[Complex_Vector_Divide.scala 44:24]
  assign io_vectorOut_7_re = io_vectorOut_7_re_divide_io_z; // @[Complex_Vector_Divide.scala 43:24]
  assign io_vectorOut_7_im = io_vectorOut_7_im_divide_io_z; // @[Complex_Vector_Divide.scala 44:24]
  assign io_vectorOut_8_re = io_vectorOut_8_re_divide_io_z; // @[Complex_Vector_Divide.scala 43:24]
  assign io_vectorOut_8_im = io_vectorOut_8_im_divide_io_z; // @[Complex_Vector_Divide.scala 44:24]
  assign io_vectorOut_9_re = io_vectorOut_9_re_divide_io_z; // @[Complex_Vector_Divide.scala 43:24]
  assign io_vectorOut_9_im = io_vectorOut_9_im_divide_io_z; // @[Complex_Vector_Divide.scala 44:24]
  assign io_vectorOut_10_re = io_vectorOut_10_re_divide_io_z; // @[Complex_Vector_Divide.scala 43:24]
  assign io_vectorOut_10_im = io_vectorOut_10_im_divide_io_z; // @[Complex_Vector_Divide.scala 44:24]
  assign io_vectorOut_11_re = io_vectorOut_11_re_divide_io_z; // @[Complex_Vector_Divide.scala 43:24]
  assign io_vectorOut_11_im = io_vectorOut_11_im_divide_io_z; // @[Complex_Vector_Divide.scala 44:24]
  assign io_vectorOut_12_re = io_vectorOut_12_re_divide_io_z; // @[Complex_Vector_Divide.scala 43:24]
  assign io_vectorOut_12_im = io_vectorOut_12_im_divide_io_z; // @[Complex_Vector_Divide.scala 44:24]
  assign io_vectorOut_13_re = io_vectorOut_13_re_divide_io_z; // @[Complex_Vector_Divide.scala 43:24]
  assign io_vectorOut_13_im = io_vectorOut_13_im_divide_io_z; // @[Complex_Vector_Divide.scala 44:24]
  assign io_vectorOut_14_re = io_vectorOut_14_re_divide_io_z; // @[Complex_Vector_Divide.scala 43:24]
  assign io_vectorOut_14_im = io_vectorOut_14_im_divide_io_z; // @[Complex_Vector_Divide.scala 44:24]
  assign io_vectorOut_15_re = io_vectorOut_15_re_divide_io_z; // @[Complex_Vector_Divide.scala 43:24]
  assign io_vectorOut_15_im = io_vectorOut_15_im_divide_io_z; // @[Complex_Vector_Divide.scala 44:24]
  assign io_vectorOut_0_re_divide_clock = clock;
  assign io_vectorOut_0_re_divide_reset = reset;
  assign io_vectorOut_0_re_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_0_re_divide_io_y = io_dividedVector_0_re; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_0_im_divide_clock = clock;
  assign io_vectorOut_0_im_divide_reset = reset;
  assign io_vectorOut_0_im_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_0_im_divide_io_y = io_dividedVector_0_im; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_1_re_divide_clock = clock;
  assign io_vectorOut_1_re_divide_reset = reset;
  assign io_vectorOut_1_re_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_1_re_divide_io_y = io_dividedVector_1_re; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_1_im_divide_clock = clock;
  assign io_vectorOut_1_im_divide_reset = reset;
  assign io_vectorOut_1_im_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_1_im_divide_io_y = io_dividedVector_1_im; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_2_re_divide_clock = clock;
  assign io_vectorOut_2_re_divide_reset = reset;
  assign io_vectorOut_2_re_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_2_re_divide_io_y = io_dividedVector_2_re; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_2_im_divide_clock = clock;
  assign io_vectorOut_2_im_divide_reset = reset;
  assign io_vectorOut_2_im_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_2_im_divide_io_y = io_dividedVector_2_im; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_3_re_divide_clock = clock;
  assign io_vectorOut_3_re_divide_reset = reset;
  assign io_vectorOut_3_re_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_3_re_divide_io_y = io_dividedVector_3_re; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_3_im_divide_clock = clock;
  assign io_vectorOut_3_im_divide_reset = reset;
  assign io_vectorOut_3_im_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_3_im_divide_io_y = io_dividedVector_3_im; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_4_re_divide_clock = clock;
  assign io_vectorOut_4_re_divide_reset = reset;
  assign io_vectorOut_4_re_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_4_re_divide_io_y = io_dividedVector_4_re; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_4_im_divide_clock = clock;
  assign io_vectorOut_4_im_divide_reset = reset;
  assign io_vectorOut_4_im_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_4_im_divide_io_y = io_dividedVector_4_im; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_5_re_divide_clock = clock;
  assign io_vectorOut_5_re_divide_reset = reset;
  assign io_vectorOut_5_re_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_5_re_divide_io_y = io_dividedVector_5_re; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_5_im_divide_clock = clock;
  assign io_vectorOut_5_im_divide_reset = reset;
  assign io_vectorOut_5_im_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_5_im_divide_io_y = io_dividedVector_5_im; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_6_re_divide_clock = clock;
  assign io_vectorOut_6_re_divide_reset = reset;
  assign io_vectorOut_6_re_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_6_re_divide_io_y = io_dividedVector_6_re; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_6_im_divide_clock = clock;
  assign io_vectorOut_6_im_divide_reset = reset;
  assign io_vectorOut_6_im_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_6_im_divide_io_y = io_dividedVector_6_im; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_7_re_divide_clock = clock;
  assign io_vectorOut_7_re_divide_reset = reset;
  assign io_vectorOut_7_re_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_7_re_divide_io_y = io_dividedVector_7_re; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_7_im_divide_clock = clock;
  assign io_vectorOut_7_im_divide_reset = reset;
  assign io_vectorOut_7_im_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_7_im_divide_io_y = io_dividedVector_7_im; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_8_re_divide_clock = clock;
  assign io_vectorOut_8_re_divide_reset = reset;
  assign io_vectorOut_8_re_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_8_re_divide_io_y = io_dividedVector_8_re; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_8_im_divide_clock = clock;
  assign io_vectorOut_8_im_divide_reset = reset;
  assign io_vectorOut_8_im_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_8_im_divide_io_y = io_dividedVector_8_im; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_9_re_divide_clock = clock;
  assign io_vectorOut_9_re_divide_reset = reset;
  assign io_vectorOut_9_re_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_9_re_divide_io_y = io_dividedVector_9_re; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_9_im_divide_clock = clock;
  assign io_vectorOut_9_im_divide_reset = reset;
  assign io_vectorOut_9_im_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_9_im_divide_io_y = io_dividedVector_9_im; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_10_re_divide_clock = clock;
  assign io_vectorOut_10_re_divide_reset = reset;
  assign io_vectorOut_10_re_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_10_re_divide_io_y = io_dividedVector_10_re; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_10_im_divide_clock = clock;
  assign io_vectorOut_10_im_divide_reset = reset;
  assign io_vectorOut_10_im_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_10_im_divide_io_y = io_dividedVector_10_im; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_11_re_divide_clock = clock;
  assign io_vectorOut_11_re_divide_reset = reset;
  assign io_vectorOut_11_re_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_11_re_divide_io_y = io_dividedVector_11_re; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_11_im_divide_clock = clock;
  assign io_vectorOut_11_im_divide_reset = reset;
  assign io_vectorOut_11_im_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_11_im_divide_io_y = io_dividedVector_11_im; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_12_re_divide_clock = clock;
  assign io_vectorOut_12_re_divide_reset = reset;
  assign io_vectorOut_12_re_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_12_re_divide_io_y = io_dividedVector_12_re; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_12_im_divide_clock = clock;
  assign io_vectorOut_12_im_divide_reset = reset;
  assign io_vectorOut_12_im_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_12_im_divide_io_y = io_dividedVector_12_im; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_13_re_divide_clock = clock;
  assign io_vectorOut_13_re_divide_reset = reset;
  assign io_vectorOut_13_re_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_13_re_divide_io_y = io_dividedVector_13_re; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_13_im_divide_clock = clock;
  assign io_vectorOut_13_im_divide_reset = reset;
  assign io_vectorOut_13_im_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_13_im_divide_io_y = io_dividedVector_13_im; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_14_re_divide_clock = clock;
  assign io_vectorOut_14_re_divide_reset = reset;
  assign io_vectorOut_14_re_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_14_re_divide_io_y = io_dividedVector_14_re; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_14_im_divide_clock = clock;
  assign io_vectorOut_14_im_divide_reset = reset;
  assign io_vectorOut_14_im_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_14_im_divide_io_y = io_dividedVector_14_im; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_15_re_divide_clock = clock;
  assign io_vectorOut_15_re_divide_reset = reset;
  assign io_vectorOut_15_re_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_15_re_divide_io_y = io_dividedVector_15_re; // @[Cordic_LV.scala 213:17]
  assign io_vectorOut_15_im_divide_clock = clock;
  assign io_vectorOut_15_im_divide_reset = reset;
  assign io_vectorOut_15_im_divide_io_x = 64'sh200000000; // @[Cordic_LV.scala 212:17]
  assign io_vectorOut_15_im_divide_io_y = io_dividedVector_15_im; // @[Cordic_LV.scala 213:17]
endmodule
module R_matirx_estimation(
  input         clock,
  input         reset,
  input         io_reset,
  input         io_ready,
  input  [63:0] io_matrixIn_0_re,
  input  [63:0] io_matrixIn_0_im,
  input  [63:0] io_matrixIn_1_re,
  input  [63:0] io_matrixIn_1_im,
  input  [63:0] io_matrixIn_2_re,
  input  [63:0] io_matrixIn_2_im,
  input  [63:0] io_matrixIn_3_re,
  input  [63:0] io_matrixIn_3_im,
  input  [63:0] io_matrixIn_4_re,
  input  [63:0] io_matrixIn_4_im,
  input  [63:0] io_matrixIn_5_re,
  input  [63:0] io_matrixIn_5_im,
  input  [63:0] io_matrixIn_6_re,
  input  [63:0] io_matrixIn_6_im,
  input  [63:0] io_matrixIn_7_re,
  input  [63:0] io_matrixIn_7_im,
  output [63:0] io_matrixOut_0_re,
  output [63:0] io_matrixOut_0_im,
  output [63:0] io_matrixOut_1_re,
  output [63:0] io_matrixOut_1_im,
  output [63:0] io_matrixOut_2_re,
  output [63:0] io_matrixOut_2_im,
  output [63:0] io_matrixOut_3_re,
  output [63:0] io_matrixOut_3_im,
  output [63:0] io_matrixOut_4_re,
  output [63:0] io_matrixOut_4_im,
  output [63:0] io_matrixOut_5_re,
  output [63:0] io_matrixOut_5_im,
  output [63:0] io_matrixOut_6_re,
  output [63:0] io_matrixOut_6_im,
  output [63:0] io_matrixOut_7_re,
  output [63:0] io_matrixOut_7_im,
  output [63:0] io_matrixOut_8_re,
  output [63:0] io_matrixOut_8_im,
  output [63:0] io_matrixOut_9_re,
  output [63:0] io_matrixOut_9_im,
  output [63:0] io_matrixOut_10_re,
  output [63:0] io_matrixOut_10_im,
  output [63:0] io_matrixOut_11_re,
  output [63:0] io_matrixOut_11_im,
  output [63:0] io_matrixOut_12_re,
  output [63:0] io_matrixOut_12_im,
  output [63:0] io_matrixOut_13_re,
  output [63:0] io_matrixOut_13_im,
  output [63:0] io_matrixOut_14_re,
  output [63:0] io_matrixOut_14_im,
  output [63:0] io_matrixOut_15_re,
  output [63:0] io_matrixOut_15_im,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
`endif // RANDOMIZE_REG_INIT
  wire  complex_matirx_mul_unit_clock; // @[R_Matrix_Estimation.scala 33:54]
  wire  complex_matirx_mul_unit_io_reset; // @[R_Matrix_Estimation.scala 33:54]
  wire  complex_matirx_mul_unit_io_ready; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_0_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_0_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_1_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_1_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_2_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_2_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_3_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_3_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixB_0_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixB_0_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixB_1_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixB_1_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixB_2_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixB_2_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixB_3_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixB_3_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_0_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_0_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_1_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_1_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_2_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_2_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_3_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_3_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_4_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_4_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_5_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_5_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_6_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_6_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_7_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_7_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_8_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_8_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_9_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_9_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_10_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_10_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_11_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_11_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_12_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_12_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_13_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_13_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_14_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_14_im; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_15_re; // @[R_Matrix_Estimation.scala 33:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_15_im; // @[R_Matrix_Estimation.scala 33:54]
  wire  complex_matirx_mul_unit_io_valid; // @[R_Matrix_Estimation.scala 33:54]
  wire  complex_vector_divide_fixedPoint_unit_clock; // @[R_Matrix_Estimation.scala 34:87]
  wire  complex_vector_divide_fixedPoint_unit_reset; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_0_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_0_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_1_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_1_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_2_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_2_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_3_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_3_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_4_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_4_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_5_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_5_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_6_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_6_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_7_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_7_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_8_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_8_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_9_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_9_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_10_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_10_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_11_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_11_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_12_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_12_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_13_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_13_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_14_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_14_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_15_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_dividedVector_15_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_0_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_0_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_1_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_1_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_2_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_2_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_3_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_3_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_4_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_4_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_5_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_5_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_6_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_6_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_7_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_7_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_8_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_8_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_9_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_9_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_10_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_10_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_11_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_11_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_12_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_12_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_13_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_13_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_14_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_14_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_15_re; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] complex_vector_divide_fixedPoint_unit_io_vectorOut_15_im; // @[R_Matrix_Estimation.scala 34:87]
  wire [63:0] matrix_mul_res_reg_0_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_0_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_0_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_0_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_0_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_0_add_io_res_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_1_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_1_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_1_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_1_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_1_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_1_add_io_res_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_2_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_2_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_2_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_2_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_2_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_2_add_io_res_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_3_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_3_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_3_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_3_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_3_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_3_add_io_res_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_4_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_4_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_4_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_4_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_4_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_4_add_io_res_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_5_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_5_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_5_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_5_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_5_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_5_add_io_res_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_6_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_6_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_6_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_6_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_6_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_6_add_io_res_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_7_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_7_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_7_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_7_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_7_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_7_add_io_res_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_8_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_8_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_8_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_8_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_8_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_8_add_io_res_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_9_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_9_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_9_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_9_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_9_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_9_add_io_res_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_10_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_10_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_10_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_10_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_10_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_10_add_io_res_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_11_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_11_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_11_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_11_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_11_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_11_add_io_res_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_12_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_12_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_12_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_12_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_12_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_12_add_io_res_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_13_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_13_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_13_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_13_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_13_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_13_add_io_res_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_14_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_14_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_14_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_14_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_14_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_14_add_io_res_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_15_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_15_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_15_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_15_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_15_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [63:0] matrix_mul_res_reg_15_add_io_res_im; // @[Complex_Operater.scala 13:21]
  reg [63:0] matrix_x_reg_0_re; // @[R_Matrix_Estimation.scala 28:39]
  reg [63:0] matrix_x_reg_0_im; // @[R_Matrix_Estimation.scala 28:39]
  reg [63:0] matrix_x_reg_1_re; // @[R_Matrix_Estimation.scala 28:39]
  reg [63:0] matrix_x_reg_1_im; // @[R_Matrix_Estimation.scala 28:39]
  reg [63:0] matrix_x_reg_2_re; // @[R_Matrix_Estimation.scala 28:39]
  reg [63:0] matrix_x_reg_2_im; // @[R_Matrix_Estimation.scala 28:39]
  reg [63:0] matrix_x_reg_3_re; // @[R_Matrix_Estimation.scala 28:39]
  reg [63:0] matrix_x_reg_3_im; // @[R_Matrix_Estimation.scala 28:39]
  reg [63:0] matrix_x_reg_4_re; // @[R_Matrix_Estimation.scala 28:39]
  reg [63:0] matrix_x_reg_4_im; // @[R_Matrix_Estimation.scala 28:39]
  reg [63:0] matrix_x_reg_5_re; // @[R_Matrix_Estimation.scala 28:39]
  reg [63:0] matrix_x_reg_5_im; // @[R_Matrix_Estimation.scala 28:39]
  reg [63:0] matrix_x_reg_6_re; // @[R_Matrix_Estimation.scala 28:39]
  reg [63:0] matrix_x_reg_6_im; // @[R_Matrix_Estimation.scala 28:39]
  reg [63:0] matrix_x_reg_7_re; // @[R_Matrix_Estimation.scala 28:39]
  reg [63:0] matrix_x_reg_7_im; // @[R_Matrix_Estimation.scala 28:39]
  reg [63:0] matrix_mul_res_reg_0_re; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_0_im; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_1_re; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_1_im; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_2_re; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_2_im; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_3_re; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_3_im; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_4_re; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_4_im; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_5_re; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_5_im; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_6_re; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_6_im; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_7_re; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_7_im; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_8_re; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_8_im; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_9_re; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_9_im; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_10_re; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_10_im; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_11_re; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_11_im; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_12_re; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_12_im; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_13_re; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_13_im; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_14_re; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_14_im; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_15_re; // @[R_Matrix_Estimation.scala 29:45]
  reg [63:0] matrix_mul_res_reg_15_im; // @[R_Matrix_Estimation.scala 29:45]
  reg [7:0] status; // @[R_Matrix_Estimation.scala 30:29]
  reg [2:0] mul_cnt; // @[R_Matrix_Estimation.scala 31:30]
  wire [4:0] _complex_matirx_mul_unit_io_matrixA_0_T = mul_cnt * 2'h2; // @[R_Matrix_Estimation.scala 62:71]
  wire [6:0] _complex_matirx_mul_unit_io_matrixA_0_T_1 = _complex_matirx_mul_unit_io_matrixA_0_T * 2'h2; // @[R_Matrix_Estimation.scala 62:77]
  wire [7:0] _complex_matirx_mul_unit_io_matrixA_0_T_2 = {{1'd0}, _complex_matirx_mul_unit_io_matrixA_0_T_1}; // @[R_Matrix_Estimation.scala 62:83]
  wire [63:0] _GEN_1 = 3'h1 == _complex_matirx_mul_unit_io_matrixA_0_T_2[2:0] ? $signed(matrix_x_reg_1_im) : $signed(
    matrix_x_reg_0_im); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_2 = 3'h2 == _complex_matirx_mul_unit_io_matrixA_0_T_2[2:0] ? $signed(matrix_x_reg_2_im) : $signed(
    _GEN_1); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_3 = 3'h3 == _complex_matirx_mul_unit_io_matrixA_0_T_2[2:0] ? $signed(matrix_x_reg_3_im) : $signed(
    _GEN_2); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_4 = 3'h4 == _complex_matirx_mul_unit_io_matrixA_0_T_2[2:0] ? $signed(matrix_x_reg_4_im) : $signed(
    _GEN_3); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_5 = 3'h5 == _complex_matirx_mul_unit_io_matrixA_0_T_2[2:0] ? $signed(matrix_x_reg_5_im) : $signed(
    _GEN_4); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_6 = 3'h6 == _complex_matirx_mul_unit_io_matrixA_0_T_2[2:0] ? $signed(matrix_x_reg_6_im) : $signed(
    _GEN_5); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_7 = 3'h7 == _complex_matirx_mul_unit_io_matrixA_0_T_2[2:0] ? $signed(matrix_x_reg_7_im) : $signed(
    _GEN_6); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_9 = 3'h1 == _complex_matirx_mul_unit_io_matrixA_0_T_2[2:0] ? $signed(matrix_x_reg_1_re) : $signed(
    matrix_x_reg_0_re); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_10 = 3'h2 == _complex_matirx_mul_unit_io_matrixA_0_T_2[2:0] ? $signed(matrix_x_reg_2_re) : $signed(
    _GEN_9); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_11 = 3'h3 == _complex_matirx_mul_unit_io_matrixA_0_T_2[2:0] ? $signed(matrix_x_reg_3_re) : $signed(
    _GEN_10); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_12 = 3'h4 == _complex_matirx_mul_unit_io_matrixA_0_T_2[2:0] ? $signed(matrix_x_reg_4_re) : $signed(
    _GEN_11); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_13 = 3'h5 == _complex_matirx_mul_unit_io_matrixA_0_T_2[2:0] ? $signed(matrix_x_reg_5_re) : $signed(
    _GEN_12); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_14 = 3'h6 == _complex_matirx_mul_unit_io_matrixA_0_T_2[2:0] ? $signed(matrix_x_reg_6_re) : $signed(
    _GEN_13); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [6:0] _complex_matirx_mul_unit_io_matrixA_1_T_3 = _complex_matirx_mul_unit_io_matrixA_0_T_1 + 7'h1; // @[R_Matrix_Estimation.scala 62:83]
  wire [63:0] _GEN_33 = 3'h1 == _complex_matirx_mul_unit_io_matrixA_1_T_3[2:0] ? $signed(matrix_x_reg_1_im) : $signed(
    matrix_x_reg_0_im); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_34 = 3'h2 == _complex_matirx_mul_unit_io_matrixA_1_T_3[2:0] ? $signed(matrix_x_reg_2_im) : $signed(
    _GEN_33); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_35 = 3'h3 == _complex_matirx_mul_unit_io_matrixA_1_T_3[2:0] ? $signed(matrix_x_reg_3_im) : $signed(
    _GEN_34); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_36 = 3'h4 == _complex_matirx_mul_unit_io_matrixA_1_T_3[2:0] ? $signed(matrix_x_reg_4_im) : $signed(
    _GEN_35); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_37 = 3'h5 == _complex_matirx_mul_unit_io_matrixA_1_T_3[2:0] ? $signed(matrix_x_reg_5_im) : $signed(
    _GEN_36); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_38 = 3'h6 == _complex_matirx_mul_unit_io_matrixA_1_T_3[2:0] ? $signed(matrix_x_reg_6_im) : $signed(
    _GEN_37); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_39 = 3'h7 == _complex_matirx_mul_unit_io_matrixA_1_T_3[2:0] ? $signed(matrix_x_reg_7_im) : $signed(
    _GEN_38); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_41 = 3'h1 == _complex_matirx_mul_unit_io_matrixA_1_T_3[2:0] ? $signed(matrix_x_reg_1_re) : $signed(
    matrix_x_reg_0_re); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_42 = 3'h2 == _complex_matirx_mul_unit_io_matrixA_1_T_3[2:0] ? $signed(matrix_x_reg_2_re) : $signed(
    _GEN_41); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_43 = 3'h3 == _complex_matirx_mul_unit_io_matrixA_1_T_3[2:0] ? $signed(matrix_x_reg_3_re) : $signed(
    _GEN_42); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_44 = 3'h4 == _complex_matirx_mul_unit_io_matrixA_1_T_3[2:0] ? $signed(matrix_x_reg_4_re) : $signed(
    _GEN_43); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_45 = 3'h5 == _complex_matirx_mul_unit_io_matrixA_1_T_3[2:0] ? $signed(matrix_x_reg_5_re) : $signed(
    _GEN_44); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_46 = 3'h6 == _complex_matirx_mul_unit_io_matrixA_1_T_3[2:0] ? $signed(matrix_x_reg_6_re) : $signed(
    _GEN_45); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [6:0] _complex_matirx_mul_unit_io_matrixA_2_T_3 = _complex_matirx_mul_unit_io_matrixA_0_T_1 + 7'h2; // @[R_Matrix_Estimation.scala 62:83]
  wire [63:0] _GEN_65 = 3'h1 == _complex_matirx_mul_unit_io_matrixA_2_T_3[2:0] ? $signed(matrix_x_reg_1_im) : $signed(
    matrix_x_reg_0_im); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_66 = 3'h2 == _complex_matirx_mul_unit_io_matrixA_2_T_3[2:0] ? $signed(matrix_x_reg_2_im) : $signed(
    _GEN_65); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_67 = 3'h3 == _complex_matirx_mul_unit_io_matrixA_2_T_3[2:0] ? $signed(matrix_x_reg_3_im) : $signed(
    _GEN_66); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_68 = 3'h4 == _complex_matirx_mul_unit_io_matrixA_2_T_3[2:0] ? $signed(matrix_x_reg_4_im) : $signed(
    _GEN_67); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_69 = 3'h5 == _complex_matirx_mul_unit_io_matrixA_2_T_3[2:0] ? $signed(matrix_x_reg_5_im) : $signed(
    _GEN_68); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_70 = 3'h6 == _complex_matirx_mul_unit_io_matrixA_2_T_3[2:0] ? $signed(matrix_x_reg_6_im) : $signed(
    _GEN_69); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_71 = 3'h7 == _complex_matirx_mul_unit_io_matrixA_2_T_3[2:0] ? $signed(matrix_x_reg_7_im) : $signed(
    _GEN_70); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_73 = 3'h1 == _complex_matirx_mul_unit_io_matrixA_2_T_3[2:0] ? $signed(matrix_x_reg_1_re) : $signed(
    matrix_x_reg_0_re); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_74 = 3'h2 == _complex_matirx_mul_unit_io_matrixA_2_T_3[2:0] ? $signed(matrix_x_reg_2_re) : $signed(
    _GEN_73); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_75 = 3'h3 == _complex_matirx_mul_unit_io_matrixA_2_T_3[2:0] ? $signed(matrix_x_reg_3_re) : $signed(
    _GEN_74); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_76 = 3'h4 == _complex_matirx_mul_unit_io_matrixA_2_T_3[2:0] ? $signed(matrix_x_reg_4_re) : $signed(
    _GEN_75); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_77 = 3'h5 == _complex_matirx_mul_unit_io_matrixA_2_T_3[2:0] ? $signed(matrix_x_reg_5_re) : $signed(
    _GEN_76); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_78 = 3'h6 == _complex_matirx_mul_unit_io_matrixA_2_T_3[2:0] ? $signed(matrix_x_reg_6_re) : $signed(
    _GEN_77); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [6:0] _complex_matirx_mul_unit_io_matrixA_3_T_3 = _complex_matirx_mul_unit_io_matrixA_0_T_1 + 7'h3; // @[R_Matrix_Estimation.scala 62:83]
  wire [63:0] _GEN_97 = 3'h1 == _complex_matirx_mul_unit_io_matrixA_3_T_3[2:0] ? $signed(matrix_x_reg_1_im) : $signed(
    matrix_x_reg_0_im); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_98 = 3'h2 == _complex_matirx_mul_unit_io_matrixA_3_T_3[2:0] ? $signed(matrix_x_reg_2_im) : $signed(
    _GEN_97); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_99 = 3'h3 == _complex_matirx_mul_unit_io_matrixA_3_T_3[2:0] ? $signed(matrix_x_reg_3_im) : $signed(
    _GEN_98); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_100 = 3'h4 == _complex_matirx_mul_unit_io_matrixA_3_T_3[2:0] ? $signed(matrix_x_reg_4_im) : $signed(
    _GEN_99); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_101 = 3'h5 == _complex_matirx_mul_unit_io_matrixA_3_T_3[2:0] ? $signed(matrix_x_reg_5_im) : $signed(
    _GEN_100); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_102 = 3'h6 == _complex_matirx_mul_unit_io_matrixA_3_T_3[2:0] ? $signed(matrix_x_reg_6_im) : $signed(
    _GEN_101); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_103 = 3'h7 == _complex_matirx_mul_unit_io_matrixA_3_T_3[2:0] ? $signed(matrix_x_reg_7_im) : $signed(
    _GEN_102); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_105 = 3'h1 == _complex_matirx_mul_unit_io_matrixA_3_T_3[2:0] ? $signed(matrix_x_reg_1_re) : $signed(
    matrix_x_reg_0_re); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_106 = 3'h2 == _complex_matirx_mul_unit_io_matrixA_3_T_3[2:0] ? $signed(matrix_x_reg_2_re) : $signed(
    _GEN_105); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_107 = 3'h3 == _complex_matirx_mul_unit_io_matrixA_3_T_3[2:0] ? $signed(matrix_x_reg_3_re) : $signed(
    _GEN_106); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_108 = 3'h4 == _complex_matirx_mul_unit_io_matrixA_3_T_3[2:0] ? $signed(matrix_x_reg_4_re) : $signed(
    _GEN_107); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_109 = 3'h5 == _complex_matirx_mul_unit_io_matrixA_3_T_3[2:0] ? $signed(matrix_x_reg_5_re) : $signed(
    _GEN_108); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [63:0] _GEN_110 = 3'h6 == _complex_matirx_mul_unit_io_matrixA_3_T_3[2:0] ? $signed(matrix_x_reg_6_re) : $signed(
    _GEN_109); // @[R_Matrix_Estimation.scala 62:{47,47}]
  wire [2:0] _mul_cnt_T_1 = mul_cnt + 3'h1; // @[R_Matrix_Estimation.scala 78:30]
  wire [1:0] _GEN_128 = mul_cnt == 3'h1 ? 2'h3 : 2'h1; // @[R_Matrix_Estimation.scala 74:37 75:18 77:18]
  wire [2:0] _GEN_129 = mul_cnt == 3'h1 ? mul_cnt : _mul_cnt_T_1; // @[R_Matrix_Estimation.scala 31:30 74:37 78:19]
  wire [63:0] _GEN_130 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_0_add_io_res_im) : $signed(
    matrix_mul_res_reg_0_im); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_131 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_0_add_io_res_re) : $signed(
    matrix_mul_res_reg_0_re); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_132 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_1_add_io_res_im) : $signed(
    matrix_mul_res_reg_1_im); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_133 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_1_add_io_res_re) : $signed(
    matrix_mul_res_reg_1_re); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_134 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_2_add_io_res_im) : $signed(
    matrix_mul_res_reg_2_im); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_135 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_2_add_io_res_re) : $signed(
    matrix_mul_res_reg_2_re); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_136 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_3_add_io_res_im) : $signed(
    matrix_mul_res_reg_3_im); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_137 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_3_add_io_res_re) : $signed(
    matrix_mul_res_reg_3_re); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_138 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_4_add_io_res_im) : $signed(
    matrix_mul_res_reg_4_im); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_139 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_4_add_io_res_re) : $signed(
    matrix_mul_res_reg_4_re); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_140 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_5_add_io_res_im) : $signed(
    matrix_mul_res_reg_5_im); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_141 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_5_add_io_res_re) : $signed(
    matrix_mul_res_reg_5_re); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_142 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_6_add_io_res_im) : $signed(
    matrix_mul_res_reg_6_im); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_143 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_6_add_io_res_re) : $signed(
    matrix_mul_res_reg_6_re); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_144 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_7_add_io_res_im) : $signed(
    matrix_mul_res_reg_7_im); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_145 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_7_add_io_res_re) : $signed(
    matrix_mul_res_reg_7_re); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_146 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_8_add_io_res_im) : $signed(
    matrix_mul_res_reg_8_im); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_147 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_8_add_io_res_re) : $signed(
    matrix_mul_res_reg_8_re); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_148 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_9_add_io_res_im) : $signed(
    matrix_mul_res_reg_9_im); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_149 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_9_add_io_res_re) : $signed(
    matrix_mul_res_reg_9_re); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_150 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_10_add_io_res_im) : $signed(
    matrix_mul_res_reg_10_im); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_151 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_10_add_io_res_re) : $signed(
    matrix_mul_res_reg_10_re); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_152 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_11_add_io_res_im) : $signed(
    matrix_mul_res_reg_11_im); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_153 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_11_add_io_res_re) : $signed(
    matrix_mul_res_reg_11_re); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_154 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_12_add_io_res_im) : $signed(
    matrix_mul_res_reg_12_im); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_155 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_12_add_io_res_re) : $signed(
    matrix_mul_res_reg_12_re); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_156 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_13_add_io_res_im) : $signed(
    matrix_mul_res_reg_13_im); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_157 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_13_add_io_res_re) : $signed(
    matrix_mul_res_reg_13_re); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_158 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_14_add_io_res_im) : $signed(
    matrix_mul_res_reg_14_im); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_159 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_14_add_io_res_re) : $signed(
    matrix_mul_res_reg_14_re); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_160 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_15_add_io_res_im) : $signed(
    matrix_mul_res_reg_15_im); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [63:0] _GEN_161 = complex_matirx_mul_unit_io_valid ? $signed(matrix_mul_res_reg_15_add_io_res_re) : $signed(
    matrix_mul_res_reg_15_re); // @[R_Matrix_Estimation.scala 70:46 72:35 29:45]
  wire [7:0] _GEN_162 = complex_matirx_mul_unit_io_valid ? {{6'd0}, _GEN_128} : status; // @[R_Matrix_Estimation.scala 30:29 70:46]
  wire [2:0] _GEN_163 = complex_matirx_mul_unit_io_valid ? _GEN_129 : mul_cnt; // @[R_Matrix_Estimation.scala 31:30 70:46]
  wire [7:0] _status_T_1 = status + 8'h1; // @[R_Matrix_Estimation.scala 85:24]
  wire [7:0] _GEN_164 = status < 8'h12 ? _status_T_1 : status; // @[R_Matrix_Estimation.scala 86:51 87:14 30:29]
  wire [7:0] _GEN_198 = status == 8'h3 ? _status_T_1 : _GEN_164; // @[R_Matrix_Estimation.scala 81:32 85:14]
  wire [7:0] _GEN_232 = status == 8'h2 ? _GEN_162 : _GEN_198; // @[R_Matrix_Estimation.scala 67:32]
  wire [2:0] _GEN_233 = status == 8'h2 ? _GEN_163 : mul_cnt; // @[R_Matrix_Estimation.scala 31:30 67:32]
  matrix_mul_v1 complex_matirx_mul_unit ( // @[R_Matrix_Estimation.scala 33:54]
    .clock(complex_matirx_mul_unit_clock),
    .io_reset(complex_matirx_mul_unit_io_reset),
    .io_ready(complex_matirx_mul_unit_io_ready),
    .io_matrixA_0_re(complex_matirx_mul_unit_io_matrixA_0_re),
    .io_matrixA_0_im(complex_matirx_mul_unit_io_matrixA_0_im),
    .io_matrixA_1_re(complex_matirx_mul_unit_io_matrixA_1_re),
    .io_matrixA_1_im(complex_matirx_mul_unit_io_matrixA_1_im),
    .io_matrixA_2_re(complex_matirx_mul_unit_io_matrixA_2_re),
    .io_matrixA_2_im(complex_matirx_mul_unit_io_matrixA_2_im),
    .io_matrixA_3_re(complex_matirx_mul_unit_io_matrixA_3_re),
    .io_matrixA_3_im(complex_matirx_mul_unit_io_matrixA_3_im),
    .io_matrixB_0_re(complex_matirx_mul_unit_io_matrixB_0_re),
    .io_matrixB_0_im(complex_matirx_mul_unit_io_matrixB_0_im),
    .io_matrixB_1_re(complex_matirx_mul_unit_io_matrixB_1_re),
    .io_matrixB_1_im(complex_matirx_mul_unit_io_matrixB_1_im),
    .io_matrixB_2_re(complex_matirx_mul_unit_io_matrixB_2_re),
    .io_matrixB_2_im(complex_matirx_mul_unit_io_matrixB_2_im),
    .io_matrixB_3_re(complex_matirx_mul_unit_io_matrixB_3_re),
    .io_matrixB_3_im(complex_matirx_mul_unit_io_matrixB_3_im),
    .io_matrixC_0_re(complex_matirx_mul_unit_io_matrixC_0_re),
    .io_matrixC_0_im(complex_matirx_mul_unit_io_matrixC_0_im),
    .io_matrixC_1_re(complex_matirx_mul_unit_io_matrixC_1_re),
    .io_matrixC_1_im(complex_matirx_mul_unit_io_matrixC_1_im),
    .io_matrixC_2_re(complex_matirx_mul_unit_io_matrixC_2_re),
    .io_matrixC_2_im(complex_matirx_mul_unit_io_matrixC_2_im),
    .io_matrixC_3_re(complex_matirx_mul_unit_io_matrixC_3_re),
    .io_matrixC_3_im(complex_matirx_mul_unit_io_matrixC_3_im),
    .io_matrixC_4_re(complex_matirx_mul_unit_io_matrixC_4_re),
    .io_matrixC_4_im(complex_matirx_mul_unit_io_matrixC_4_im),
    .io_matrixC_5_re(complex_matirx_mul_unit_io_matrixC_5_re),
    .io_matrixC_5_im(complex_matirx_mul_unit_io_matrixC_5_im),
    .io_matrixC_6_re(complex_matirx_mul_unit_io_matrixC_6_re),
    .io_matrixC_6_im(complex_matirx_mul_unit_io_matrixC_6_im),
    .io_matrixC_7_re(complex_matirx_mul_unit_io_matrixC_7_re),
    .io_matrixC_7_im(complex_matirx_mul_unit_io_matrixC_7_im),
    .io_matrixC_8_re(complex_matirx_mul_unit_io_matrixC_8_re),
    .io_matrixC_8_im(complex_matirx_mul_unit_io_matrixC_8_im),
    .io_matrixC_9_re(complex_matirx_mul_unit_io_matrixC_9_re),
    .io_matrixC_9_im(complex_matirx_mul_unit_io_matrixC_9_im),
    .io_matrixC_10_re(complex_matirx_mul_unit_io_matrixC_10_re),
    .io_matrixC_10_im(complex_matirx_mul_unit_io_matrixC_10_im),
    .io_matrixC_11_re(complex_matirx_mul_unit_io_matrixC_11_re),
    .io_matrixC_11_im(complex_matirx_mul_unit_io_matrixC_11_im),
    .io_matrixC_12_re(complex_matirx_mul_unit_io_matrixC_12_re),
    .io_matrixC_12_im(complex_matirx_mul_unit_io_matrixC_12_im),
    .io_matrixC_13_re(complex_matirx_mul_unit_io_matrixC_13_re),
    .io_matrixC_13_im(complex_matirx_mul_unit_io_matrixC_13_im),
    .io_matrixC_14_re(complex_matirx_mul_unit_io_matrixC_14_re),
    .io_matrixC_14_im(complex_matirx_mul_unit_io_matrixC_14_im),
    .io_matrixC_15_re(complex_matirx_mul_unit_io_matrixC_15_re),
    .io_matrixC_15_im(complex_matirx_mul_unit_io_matrixC_15_im),
    .io_valid(complex_matirx_mul_unit_io_valid)
  );
  complex_vector_divide_fixedPoint complex_vector_divide_fixedPoint_unit ( // @[R_Matrix_Estimation.scala 34:87]
    .clock(complex_vector_divide_fixedPoint_unit_clock),
    .reset(complex_vector_divide_fixedPoint_unit_reset),
    .io_dividedVector_0_re(complex_vector_divide_fixedPoint_unit_io_dividedVector_0_re),
    .io_dividedVector_0_im(complex_vector_divide_fixedPoint_unit_io_dividedVector_0_im),
    .io_dividedVector_1_re(complex_vector_divide_fixedPoint_unit_io_dividedVector_1_re),
    .io_dividedVector_1_im(complex_vector_divide_fixedPoint_unit_io_dividedVector_1_im),
    .io_dividedVector_2_re(complex_vector_divide_fixedPoint_unit_io_dividedVector_2_re),
    .io_dividedVector_2_im(complex_vector_divide_fixedPoint_unit_io_dividedVector_2_im),
    .io_dividedVector_3_re(complex_vector_divide_fixedPoint_unit_io_dividedVector_3_re),
    .io_dividedVector_3_im(complex_vector_divide_fixedPoint_unit_io_dividedVector_3_im),
    .io_dividedVector_4_re(complex_vector_divide_fixedPoint_unit_io_dividedVector_4_re),
    .io_dividedVector_4_im(complex_vector_divide_fixedPoint_unit_io_dividedVector_4_im),
    .io_dividedVector_5_re(complex_vector_divide_fixedPoint_unit_io_dividedVector_5_re),
    .io_dividedVector_5_im(complex_vector_divide_fixedPoint_unit_io_dividedVector_5_im),
    .io_dividedVector_6_re(complex_vector_divide_fixedPoint_unit_io_dividedVector_6_re),
    .io_dividedVector_6_im(complex_vector_divide_fixedPoint_unit_io_dividedVector_6_im),
    .io_dividedVector_7_re(complex_vector_divide_fixedPoint_unit_io_dividedVector_7_re),
    .io_dividedVector_7_im(complex_vector_divide_fixedPoint_unit_io_dividedVector_7_im),
    .io_dividedVector_8_re(complex_vector_divide_fixedPoint_unit_io_dividedVector_8_re),
    .io_dividedVector_8_im(complex_vector_divide_fixedPoint_unit_io_dividedVector_8_im),
    .io_dividedVector_9_re(complex_vector_divide_fixedPoint_unit_io_dividedVector_9_re),
    .io_dividedVector_9_im(complex_vector_divide_fixedPoint_unit_io_dividedVector_9_im),
    .io_dividedVector_10_re(complex_vector_divide_fixedPoint_unit_io_dividedVector_10_re),
    .io_dividedVector_10_im(complex_vector_divide_fixedPoint_unit_io_dividedVector_10_im),
    .io_dividedVector_11_re(complex_vector_divide_fixedPoint_unit_io_dividedVector_11_re),
    .io_dividedVector_11_im(complex_vector_divide_fixedPoint_unit_io_dividedVector_11_im),
    .io_dividedVector_12_re(complex_vector_divide_fixedPoint_unit_io_dividedVector_12_re),
    .io_dividedVector_12_im(complex_vector_divide_fixedPoint_unit_io_dividedVector_12_im),
    .io_dividedVector_13_re(complex_vector_divide_fixedPoint_unit_io_dividedVector_13_re),
    .io_dividedVector_13_im(complex_vector_divide_fixedPoint_unit_io_dividedVector_13_im),
    .io_dividedVector_14_re(complex_vector_divide_fixedPoint_unit_io_dividedVector_14_re),
    .io_dividedVector_14_im(complex_vector_divide_fixedPoint_unit_io_dividedVector_14_im),
    .io_dividedVector_15_re(complex_vector_divide_fixedPoint_unit_io_dividedVector_15_re),
    .io_dividedVector_15_im(complex_vector_divide_fixedPoint_unit_io_dividedVector_15_im),
    .io_vectorOut_0_re(complex_vector_divide_fixedPoint_unit_io_vectorOut_0_re),
    .io_vectorOut_0_im(complex_vector_divide_fixedPoint_unit_io_vectorOut_0_im),
    .io_vectorOut_1_re(complex_vector_divide_fixedPoint_unit_io_vectorOut_1_re),
    .io_vectorOut_1_im(complex_vector_divide_fixedPoint_unit_io_vectorOut_1_im),
    .io_vectorOut_2_re(complex_vector_divide_fixedPoint_unit_io_vectorOut_2_re),
    .io_vectorOut_2_im(complex_vector_divide_fixedPoint_unit_io_vectorOut_2_im),
    .io_vectorOut_3_re(complex_vector_divide_fixedPoint_unit_io_vectorOut_3_re),
    .io_vectorOut_3_im(complex_vector_divide_fixedPoint_unit_io_vectorOut_3_im),
    .io_vectorOut_4_re(complex_vector_divide_fixedPoint_unit_io_vectorOut_4_re),
    .io_vectorOut_4_im(complex_vector_divide_fixedPoint_unit_io_vectorOut_4_im),
    .io_vectorOut_5_re(complex_vector_divide_fixedPoint_unit_io_vectorOut_5_re),
    .io_vectorOut_5_im(complex_vector_divide_fixedPoint_unit_io_vectorOut_5_im),
    .io_vectorOut_6_re(complex_vector_divide_fixedPoint_unit_io_vectorOut_6_re),
    .io_vectorOut_6_im(complex_vector_divide_fixedPoint_unit_io_vectorOut_6_im),
    .io_vectorOut_7_re(complex_vector_divide_fixedPoint_unit_io_vectorOut_7_re),
    .io_vectorOut_7_im(complex_vector_divide_fixedPoint_unit_io_vectorOut_7_im),
    .io_vectorOut_8_re(complex_vector_divide_fixedPoint_unit_io_vectorOut_8_re),
    .io_vectorOut_8_im(complex_vector_divide_fixedPoint_unit_io_vectorOut_8_im),
    .io_vectorOut_9_re(complex_vector_divide_fixedPoint_unit_io_vectorOut_9_re),
    .io_vectorOut_9_im(complex_vector_divide_fixedPoint_unit_io_vectorOut_9_im),
    .io_vectorOut_10_re(complex_vector_divide_fixedPoint_unit_io_vectorOut_10_re),
    .io_vectorOut_10_im(complex_vector_divide_fixedPoint_unit_io_vectorOut_10_im),
    .io_vectorOut_11_re(complex_vector_divide_fixedPoint_unit_io_vectorOut_11_re),
    .io_vectorOut_11_im(complex_vector_divide_fixedPoint_unit_io_vectorOut_11_im),
    .io_vectorOut_12_re(complex_vector_divide_fixedPoint_unit_io_vectorOut_12_re),
    .io_vectorOut_12_im(complex_vector_divide_fixedPoint_unit_io_vectorOut_12_im),
    .io_vectorOut_13_re(complex_vector_divide_fixedPoint_unit_io_vectorOut_13_re),
    .io_vectorOut_13_im(complex_vector_divide_fixedPoint_unit_io_vectorOut_13_im),
    .io_vectorOut_14_re(complex_vector_divide_fixedPoint_unit_io_vectorOut_14_re),
    .io_vectorOut_14_im(complex_vector_divide_fixedPoint_unit_io_vectorOut_14_im),
    .io_vectorOut_15_re(complex_vector_divide_fixedPoint_unit_io_vectorOut_15_re),
    .io_vectorOut_15_im(complex_vector_divide_fixedPoint_unit_io_vectorOut_15_im)
  );
  ComplexAdd matrix_mul_res_reg_0_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(matrix_mul_res_reg_0_add_io_op1_re),
    .io_op1_im(matrix_mul_res_reg_0_add_io_op1_im),
    .io_op2_re(matrix_mul_res_reg_0_add_io_op2_re),
    .io_op2_im(matrix_mul_res_reg_0_add_io_op2_im),
    .io_res_re(matrix_mul_res_reg_0_add_io_res_re),
    .io_res_im(matrix_mul_res_reg_0_add_io_res_im)
  );
  ComplexAdd matrix_mul_res_reg_1_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(matrix_mul_res_reg_1_add_io_op1_re),
    .io_op1_im(matrix_mul_res_reg_1_add_io_op1_im),
    .io_op2_re(matrix_mul_res_reg_1_add_io_op2_re),
    .io_op2_im(matrix_mul_res_reg_1_add_io_op2_im),
    .io_res_re(matrix_mul_res_reg_1_add_io_res_re),
    .io_res_im(matrix_mul_res_reg_1_add_io_res_im)
  );
  ComplexAdd matrix_mul_res_reg_2_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(matrix_mul_res_reg_2_add_io_op1_re),
    .io_op1_im(matrix_mul_res_reg_2_add_io_op1_im),
    .io_op2_re(matrix_mul_res_reg_2_add_io_op2_re),
    .io_op2_im(matrix_mul_res_reg_2_add_io_op2_im),
    .io_res_re(matrix_mul_res_reg_2_add_io_res_re),
    .io_res_im(matrix_mul_res_reg_2_add_io_res_im)
  );
  ComplexAdd matrix_mul_res_reg_3_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(matrix_mul_res_reg_3_add_io_op1_re),
    .io_op1_im(matrix_mul_res_reg_3_add_io_op1_im),
    .io_op2_re(matrix_mul_res_reg_3_add_io_op2_re),
    .io_op2_im(matrix_mul_res_reg_3_add_io_op2_im),
    .io_res_re(matrix_mul_res_reg_3_add_io_res_re),
    .io_res_im(matrix_mul_res_reg_3_add_io_res_im)
  );
  ComplexAdd matrix_mul_res_reg_4_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(matrix_mul_res_reg_4_add_io_op1_re),
    .io_op1_im(matrix_mul_res_reg_4_add_io_op1_im),
    .io_op2_re(matrix_mul_res_reg_4_add_io_op2_re),
    .io_op2_im(matrix_mul_res_reg_4_add_io_op2_im),
    .io_res_re(matrix_mul_res_reg_4_add_io_res_re),
    .io_res_im(matrix_mul_res_reg_4_add_io_res_im)
  );
  ComplexAdd matrix_mul_res_reg_5_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(matrix_mul_res_reg_5_add_io_op1_re),
    .io_op1_im(matrix_mul_res_reg_5_add_io_op1_im),
    .io_op2_re(matrix_mul_res_reg_5_add_io_op2_re),
    .io_op2_im(matrix_mul_res_reg_5_add_io_op2_im),
    .io_res_re(matrix_mul_res_reg_5_add_io_res_re),
    .io_res_im(matrix_mul_res_reg_5_add_io_res_im)
  );
  ComplexAdd matrix_mul_res_reg_6_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(matrix_mul_res_reg_6_add_io_op1_re),
    .io_op1_im(matrix_mul_res_reg_6_add_io_op1_im),
    .io_op2_re(matrix_mul_res_reg_6_add_io_op2_re),
    .io_op2_im(matrix_mul_res_reg_6_add_io_op2_im),
    .io_res_re(matrix_mul_res_reg_6_add_io_res_re),
    .io_res_im(matrix_mul_res_reg_6_add_io_res_im)
  );
  ComplexAdd matrix_mul_res_reg_7_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(matrix_mul_res_reg_7_add_io_op1_re),
    .io_op1_im(matrix_mul_res_reg_7_add_io_op1_im),
    .io_op2_re(matrix_mul_res_reg_7_add_io_op2_re),
    .io_op2_im(matrix_mul_res_reg_7_add_io_op2_im),
    .io_res_re(matrix_mul_res_reg_7_add_io_res_re),
    .io_res_im(matrix_mul_res_reg_7_add_io_res_im)
  );
  ComplexAdd matrix_mul_res_reg_8_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(matrix_mul_res_reg_8_add_io_op1_re),
    .io_op1_im(matrix_mul_res_reg_8_add_io_op1_im),
    .io_op2_re(matrix_mul_res_reg_8_add_io_op2_re),
    .io_op2_im(matrix_mul_res_reg_8_add_io_op2_im),
    .io_res_re(matrix_mul_res_reg_8_add_io_res_re),
    .io_res_im(matrix_mul_res_reg_8_add_io_res_im)
  );
  ComplexAdd matrix_mul_res_reg_9_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(matrix_mul_res_reg_9_add_io_op1_re),
    .io_op1_im(matrix_mul_res_reg_9_add_io_op1_im),
    .io_op2_re(matrix_mul_res_reg_9_add_io_op2_re),
    .io_op2_im(matrix_mul_res_reg_9_add_io_op2_im),
    .io_res_re(matrix_mul_res_reg_9_add_io_res_re),
    .io_res_im(matrix_mul_res_reg_9_add_io_res_im)
  );
  ComplexAdd matrix_mul_res_reg_10_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(matrix_mul_res_reg_10_add_io_op1_re),
    .io_op1_im(matrix_mul_res_reg_10_add_io_op1_im),
    .io_op2_re(matrix_mul_res_reg_10_add_io_op2_re),
    .io_op2_im(matrix_mul_res_reg_10_add_io_op2_im),
    .io_res_re(matrix_mul_res_reg_10_add_io_res_re),
    .io_res_im(matrix_mul_res_reg_10_add_io_res_im)
  );
  ComplexAdd matrix_mul_res_reg_11_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(matrix_mul_res_reg_11_add_io_op1_re),
    .io_op1_im(matrix_mul_res_reg_11_add_io_op1_im),
    .io_op2_re(matrix_mul_res_reg_11_add_io_op2_re),
    .io_op2_im(matrix_mul_res_reg_11_add_io_op2_im),
    .io_res_re(matrix_mul_res_reg_11_add_io_res_re),
    .io_res_im(matrix_mul_res_reg_11_add_io_res_im)
  );
  ComplexAdd matrix_mul_res_reg_12_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(matrix_mul_res_reg_12_add_io_op1_re),
    .io_op1_im(matrix_mul_res_reg_12_add_io_op1_im),
    .io_op2_re(matrix_mul_res_reg_12_add_io_op2_re),
    .io_op2_im(matrix_mul_res_reg_12_add_io_op2_im),
    .io_res_re(matrix_mul_res_reg_12_add_io_res_re),
    .io_res_im(matrix_mul_res_reg_12_add_io_res_im)
  );
  ComplexAdd matrix_mul_res_reg_13_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(matrix_mul_res_reg_13_add_io_op1_re),
    .io_op1_im(matrix_mul_res_reg_13_add_io_op1_im),
    .io_op2_re(matrix_mul_res_reg_13_add_io_op2_re),
    .io_op2_im(matrix_mul_res_reg_13_add_io_op2_im),
    .io_res_re(matrix_mul_res_reg_13_add_io_res_re),
    .io_res_im(matrix_mul_res_reg_13_add_io_res_im)
  );
  ComplexAdd matrix_mul_res_reg_14_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(matrix_mul_res_reg_14_add_io_op1_re),
    .io_op1_im(matrix_mul_res_reg_14_add_io_op1_im),
    .io_op2_re(matrix_mul_res_reg_14_add_io_op2_re),
    .io_op2_im(matrix_mul_res_reg_14_add_io_op2_im),
    .io_res_re(matrix_mul_res_reg_14_add_io_res_re),
    .io_res_im(matrix_mul_res_reg_14_add_io_res_im)
  );
  ComplexAdd matrix_mul_res_reg_15_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(matrix_mul_res_reg_15_add_io_op1_re),
    .io_op1_im(matrix_mul_res_reg_15_add_io_op1_im),
    .io_op2_re(matrix_mul_res_reg_15_add_io_op2_re),
    .io_op2_im(matrix_mul_res_reg_15_add_io_op2_im),
    .io_res_re(matrix_mul_res_reg_15_add_io_res_re),
    .io_res_im(matrix_mul_res_reg_15_add_io_res_im)
  );
  assign io_matrixOut_0_re = complex_vector_divide_fixedPoint_unit_io_vectorOut_0_re; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_0_im = complex_vector_divide_fixedPoint_unit_io_vectorOut_0_im; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_1_re = complex_vector_divide_fixedPoint_unit_io_vectorOut_1_re; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_1_im = complex_vector_divide_fixedPoint_unit_io_vectorOut_1_im; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_2_re = complex_vector_divide_fixedPoint_unit_io_vectorOut_2_re; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_2_im = complex_vector_divide_fixedPoint_unit_io_vectorOut_2_im; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_3_re = complex_vector_divide_fixedPoint_unit_io_vectorOut_3_re; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_3_im = complex_vector_divide_fixedPoint_unit_io_vectorOut_3_im; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_4_re = complex_vector_divide_fixedPoint_unit_io_vectorOut_4_re; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_4_im = complex_vector_divide_fixedPoint_unit_io_vectorOut_4_im; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_5_re = complex_vector_divide_fixedPoint_unit_io_vectorOut_5_re; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_5_im = complex_vector_divide_fixedPoint_unit_io_vectorOut_5_im; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_6_re = complex_vector_divide_fixedPoint_unit_io_vectorOut_6_re; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_6_im = complex_vector_divide_fixedPoint_unit_io_vectorOut_6_im; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_7_re = complex_vector_divide_fixedPoint_unit_io_vectorOut_7_re; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_7_im = complex_vector_divide_fixedPoint_unit_io_vectorOut_7_im; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_8_re = complex_vector_divide_fixedPoint_unit_io_vectorOut_8_re; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_8_im = complex_vector_divide_fixedPoint_unit_io_vectorOut_8_im; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_9_re = complex_vector_divide_fixedPoint_unit_io_vectorOut_9_re; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_9_im = complex_vector_divide_fixedPoint_unit_io_vectorOut_9_im; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_10_re = complex_vector_divide_fixedPoint_unit_io_vectorOut_10_re; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_10_im = complex_vector_divide_fixedPoint_unit_io_vectorOut_10_im; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_11_re = complex_vector_divide_fixedPoint_unit_io_vectorOut_11_re; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_11_im = complex_vector_divide_fixedPoint_unit_io_vectorOut_11_im; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_12_re = complex_vector_divide_fixedPoint_unit_io_vectorOut_12_re; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_12_im = complex_vector_divide_fixedPoint_unit_io_vectorOut_12_im; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_13_re = complex_vector_divide_fixedPoint_unit_io_vectorOut_13_re; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_13_im = complex_vector_divide_fixedPoint_unit_io_vectorOut_13_im; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_14_re = complex_vector_divide_fixedPoint_unit_io_vectorOut_14_re; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_14_im = complex_vector_divide_fixedPoint_unit_io_vectorOut_14_im; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_15_re = complex_vector_divide_fixedPoint_unit_io_vectorOut_15_re; // @[R_Matrix_Estimation.scala 96:16]
  assign io_matrixOut_15_im = complex_vector_divide_fixedPoint_unit_io_vectorOut_15_im; // @[R_Matrix_Estimation.scala 96:16]
  assign io_valid = status >= 8'h12; // @[R_Matrix_Estimation.scala 91:15]
  assign complex_matirx_mul_unit_clock = clock;
  assign complex_matirx_mul_unit_io_reset = io_reset; // @[R_Matrix_Estimation.scala 35:36]
  assign complex_matirx_mul_unit_io_ready = status == 8'h1; // @[R_Matrix_Estimation.scala 58:17]
  assign complex_matirx_mul_unit_io_matrixA_0_re = 3'h7 == _complex_matirx_mul_unit_io_matrixA_0_T_2[2:0] ? $signed(
    matrix_x_reg_7_re) : $signed(_GEN_14); // @[R_Matrix_Estimation.scala 62:{47,47}]
  assign complex_matirx_mul_unit_io_matrixA_0_im = 3'h7 == _complex_matirx_mul_unit_io_matrixA_0_T_2[2:0] ? $signed(
    matrix_x_reg_7_im) : $signed(_GEN_6); // @[R_Matrix_Estimation.scala 62:{47,47}]
  assign complex_matirx_mul_unit_io_matrixA_1_re = 3'h7 == _complex_matirx_mul_unit_io_matrixA_1_T_3[2:0] ? $signed(
    matrix_x_reg_7_re) : $signed(_GEN_46); // @[R_Matrix_Estimation.scala 62:{47,47}]
  assign complex_matirx_mul_unit_io_matrixA_1_im = 3'h7 == _complex_matirx_mul_unit_io_matrixA_1_T_3[2:0] ? $signed(
    matrix_x_reg_7_im) : $signed(_GEN_38); // @[R_Matrix_Estimation.scala 62:{47,47}]
  assign complex_matirx_mul_unit_io_matrixA_2_re = 3'h7 == _complex_matirx_mul_unit_io_matrixA_2_T_3[2:0] ? $signed(
    matrix_x_reg_7_re) : $signed(_GEN_78); // @[R_Matrix_Estimation.scala 62:{47,47}]
  assign complex_matirx_mul_unit_io_matrixA_2_im = 3'h7 == _complex_matirx_mul_unit_io_matrixA_2_T_3[2:0] ? $signed(
    matrix_x_reg_7_im) : $signed(_GEN_70); // @[R_Matrix_Estimation.scala 62:{47,47}]
  assign complex_matirx_mul_unit_io_matrixA_3_re = 3'h7 == _complex_matirx_mul_unit_io_matrixA_3_T_3[2:0] ? $signed(
    matrix_x_reg_7_re) : $signed(_GEN_110); // @[R_Matrix_Estimation.scala 62:{47,47}]
  assign complex_matirx_mul_unit_io_matrixA_3_im = 3'h7 == _complex_matirx_mul_unit_io_matrixA_3_T_3[2:0] ? $signed(
    matrix_x_reg_7_im) : $signed(_GEN_102); // @[R_Matrix_Estimation.scala 62:{47,47}]
  assign complex_matirx_mul_unit_io_matrixB_0_re = 3'h7 == _complex_matirx_mul_unit_io_matrixA_0_T_2[2:0] ? $signed(
    matrix_x_reg_7_re) : $signed(_GEN_14); // @[R_Matrix_Estimation.scala 63:{50,50}]
  assign complex_matirx_mul_unit_io_matrixB_0_im = 64'sh0 - $signed(_GEN_7); // @[R_Matrix_Estimation.scala 64:53]
  assign complex_matirx_mul_unit_io_matrixB_1_re = 3'h7 == _complex_matirx_mul_unit_io_matrixA_1_T_3[2:0] ? $signed(
    matrix_x_reg_7_re) : $signed(_GEN_46); // @[R_Matrix_Estimation.scala 63:{50,50}]
  assign complex_matirx_mul_unit_io_matrixB_1_im = 64'sh0 - $signed(_GEN_39); // @[R_Matrix_Estimation.scala 64:53]
  assign complex_matirx_mul_unit_io_matrixB_2_re = 3'h7 == _complex_matirx_mul_unit_io_matrixA_2_T_3[2:0] ? $signed(
    matrix_x_reg_7_re) : $signed(_GEN_78); // @[R_Matrix_Estimation.scala 63:{50,50}]
  assign complex_matirx_mul_unit_io_matrixB_2_im = 64'sh0 - $signed(_GEN_71); // @[R_Matrix_Estimation.scala 64:53]
  assign complex_matirx_mul_unit_io_matrixB_3_re = 3'h7 == _complex_matirx_mul_unit_io_matrixA_3_T_3[2:0] ? $signed(
    matrix_x_reg_7_re) : $signed(_GEN_110); // @[R_Matrix_Estimation.scala 63:{50,50}]
  assign complex_matirx_mul_unit_io_matrixB_3_im = 64'sh0 - $signed(_GEN_103); // @[R_Matrix_Estimation.scala 64:53]
  assign complex_vector_divide_fixedPoint_unit_clock = clock;
  assign complex_vector_divide_fixedPoint_unit_reset = reset;
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_0_re = matrix_mul_res_reg_0_re; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_0_im = matrix_mul_res_reg_0_im; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_1_re = matrix_mul_res_reg_1_re; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_1_im = matrix_mul_res_reg_1_im; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_2_re = matrix_mul_res_reg_2_re; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_2_im = matrix_mul_res_reg_2_im; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_3_re = matrix_mul_res_reg_3_re; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_3_im = matrix_mul_res_reg_3_im; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_4_re = matrix_mul_res_reg_4_re; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_4_im = matrix_mul_res_reg_4_im; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_5_re = matrix_mul_res_reg_5_re; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_5_im = matrix_mul_res_reg_5_im; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_6_re = matrix_mul_res_reg_6_re; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_6_im = matrix_mul_res_reg_6_im; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_7_re = matrix_mul_res_reg_7_re; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_7_im = matrix_mul_res_reg_7_im; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_8_re = matrix_mul_res_reg_8_re; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_8_im = matrix_mul_res_reg_8_im; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_9_re = matrix_mul_res_reg_9_re; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_9_im = matrix_mul_res_reg_9_im; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_10_re = matrix_mul_res_reg_10_re; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_10_im = matrix_mul_res_reg_10_im; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_11_re = matrix_mul_res_reg_11_re; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_11_im = matrix_mul_res_reg_11_im; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_12_re = matrix_mul_res_reg_12_re; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_12_im = matrix_mul_res_reg_12_im; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_13_re = matrix_mul_res_reg_13_re; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_13_im = matrix_mul_res_reg_13_im; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_14_re = matrix_mul_res_reg_14_re; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_14_im = matrix_mul_res_reg_14_im; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_15_re = matrix_mul_res_reg_15_re; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign complex_vector_divide_fixedPoint_unit_io_dividedVector_15_im = matrix_mul_res_reg_15_im; // @[R_Matrix_Estimation.scala 81:32 83:62]
  assign matrix_mul_res_reg_0_add_io_op1_re = matrix_mul_res_reg_0_re; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_0_add_io_op1_im = matrix_mul_res_reg_0_im; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_0_add_io_op2_re = complex_matirx_mul_unit_io_matrixC_0_re; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_0_add_io_op2_im = complex_matirx_mul_unit_io_matrixC_0_im; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_1_add_io_op1_re = matrix_mul_res_reg_1_re; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_1_add_io_op1_im = matrix_mul_res_reg_1_im; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_1_add_io_op2_re = complex_matirx_mul_unit_io_matrixC_1_re; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_1_add_io_op2_im = complex_matirx_mul_unit_io_matrixC_1_im; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_2_add_io_op1_re = matrix_mul_res_reg_2_re; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_2_add_io_op1_im = matrix_mul_res_reg_2_im; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_2_add_io_op2_re = complex_matirx_mul_unit_io_matrixC_2_re; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_2_add_io_op2_im = complex_matirx_mul_unit_io_matrixC_2_im; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_3_add_io_op1_re = matrix_mul_res_reg_3_re; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_3_add_io_op1_im = matrix_mul_res_reg_3_im; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_3_add_io_op2_re = complex_matirx_mul_unit_io_matrixC_3_re; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_3_add_io_op2_im = complex_matirx_mul_unit_io_matrixC_3_im; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_4_add_io_op1_re = matrix_mul_res_reg_4_re; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_4_add_io_op1_im = matrix_mul_res_reg_4_im; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_4_add_io_op2_re = complex_matirx_mul_unit_io_matrixC_4_re; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_4_add_io_op2_im = complex_matirx_mul_unit_io_matrixC_4_im; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_5_add_io_op1_re = matrix_mul_res_reg_5_re; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_5_add_io_op1_im = matrix_mul_res_reg_5_im; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_5_add_io_op2_re = complex_matirx_mul_unit_io_matrixC_5_re; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_5_add_io_op2_im = complex_matirx_mul_unit_io_matrixC_5_im; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_6_add_io_op1_re = matrix_mul_res_reg_6_re; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_6_add_io_op1_im = matrix_mul_res_reg_6_im; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_6_add_io_op2_re = complex_matirx_mul_unit_io_matrixC_6_re; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_6_add_io_op2_im = complex_matirx_mul_unit_io_matrixC_6_im; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_7_add_io_op1_re = matrix_mul_res_reg_7_re; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_7_add_io_op1_im = matrix_mul_res_reg_7_im; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_7_add_io_op2_re = complex_matirx_mul_unit_io_matrixC_7_re; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_7_add_io_op2_im = complex_matirx_mul_unit_io_matrixC_7_im; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_8_add_io_op1_re = matrix_mul_res_reg_8_re; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_8_add_io_op1_im = matrix_mul_res_reg_8_im; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_8_add_io_op2_re = complex_matirx_mul_unit_io_matrixC_8_re; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_8_add_io_op2_im = complex_matirx_mul_unit_io_matrixC_8_im; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_9_add_io_op1_re = matrix_mul_res_reg_9_re; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_9_add_io_op1_im = matrix_mul_res_reg_9_im; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_9_add_io_op2_re = complex_matirx_mul_unit_io_matrixC_9_re; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_9_add_io_op2_im = complex_matirx_mul_unit_io_matrixC_9_im; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_10_add_io_op1_re = matrix_mul_res_reg_10_re; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_10_add_io_op1_im = matrix_mul_res_reg_10_im; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_10_add_io_op2_re = complex_matirx_mul_unit_io_matrixC_10_re; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_10_add_io_op2_im = complex_matirx_mul_unit_io_matrixC_10_im; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_11_add_io_op1_re = matrix_mul_res_reg_11_re; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_11_add_io_op1_im = matrix_mul_res_reg_11_im; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_11_add_io_op2_re = complex_matirx_mul_unit_io_matrixC_11_re; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_11_add_io_op2_im = complex_matirx_mul_unit_io_matrixC_11_im; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_12_add_io_op1_re = matrix_mul_res_reg_12_re; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_12_add_io_op1_im = matrix_mul_res_reg_12_im; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_12_add_io_op2_re = complex_matirx_mul_unit_io_matrixC_12_re; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_12_add_io_op2_im = complex_matirx_mul_unit_io_matrixC_12_im; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_13_add_io_op1_re = matrix_mul_res_reg_13_re; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_13_add_io_op1_im = matrix_mul_res_reg_13_im; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_13_add_io_op2_re = complex_matirx_mul_unit_io_matrixC_13_re; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_13_add_io_op2_im = complex_matirx_mul_unit_io_matrixC_13_im; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_14_add_io_op1_re = matrix_mul_res_reg_14_re; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_14_add_io_op1_im = matrix_mul_res_reg_14_im; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_14_add_io_op2_re = complex_matirx_mul_unit_io_matrixC_14_re; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_14_add_io_op2_im = complex_matirx_mul_unit_io_matrixC_14_im; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_15_add_io_op1_re = matrix_mul_res_reg_15_re; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_15_add_io_op1_im = matrix_mul_res_reg_15_im; // @[Complex_Operater.scala 14:16]
  assign matrix_mul_res_reg_15_add_io_op2_re = complex_matirx_mul_unit_io_matrixC_15_re; // @[Complex_Operater.scala 15:16]
  assign matrix_mul_res_reg_15_add_io_op2_im = complex_matirx_mul_unit_io_matrixC_15_im; // @[Complex_Operater.scala 15:16]
  always @(posedge clock) begin
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_x_reg_0_re <= 64'sh0; // @[R_Matrix_Estimation.scala 44:26]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      matrix_x_reg_0_re <= io_matrixIn_0_re; // @[R_Matrix_Estimation.scala 54:18]
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_x_reg_0_im <= 64'sh0; // @[R_Matrix_Estimation.scala 45:26]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      matrix_x_reg_0_im <= io_matrixIn_0_im; // @[R_Matrix_Estimation.scala 54:18]
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_x_reg_1_re <= 64'sh0; // @[R_Matrix_Estimation.scala 44:26]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      matrix_x_reg_1_re <= io_matrixIn_1_re; // @[R_Matrix_Estimation.scala 54:18]
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_x_reg_1_im <= 64'sh0; // @[R_Matrix_Estimation.scala 45:26]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      matrix_x_reg_1_im <= io_matrixIn_1_im; // @[R_Matrix_Estimation.scala 54:18]
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_x_reg_2_re <= 64'sh0; // @[R_Matrix_Estimation.scala 44:26]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      matrix_x_reg_2_re <= io_matrixIn_2_re; // @[R_Matrix_Estimation.scala 54:18]
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_x_reg_2_im <= 64'sh0; // @[R_Matrix_Estimation.scala 45:26]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      matrix_x_reg_2_im <= io_matrixIn_2_im; // @[R_Matrix_Estimation.scala 54:18]
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_x_reg_3_re <= 64'sh0; // @[R_Matrix_Estimation.scala 44:26]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      matrix_x_reg_3_re <= io_matrixIn_3_re; // @[R_Matrix_Estimation.scala 54:18]
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_x_reg_3_im <= 64'sh0; // @[R_Matrix_Estimation.scala 45:26]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      matrix_x_reg_3_im <= io_matrixIn_3_im; // @[R_Matrix_Estimation.scala 54:18]
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_x_reg_4_re <= 64'sh0; // @[R_Matrix_Estimation.scala 44:26]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      matrix_x_reg_4_re <= io_matrixIn_4_re; // @[R_Matrix_Estimation.scala 54:18]
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_x_reg_4_im <= 64'sh0; // @[R_Matrix_Estimation.scala 45:26]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      matrix_x_reg_4_im <= io_matrixIn_4_im; // @[R_Matrix_Estimation.scala 54:18]
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_x_reg_5_re <= 64'sh0; // @[R_Matrix_Estimation.scala 44:26]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      matrix_x_reg_5_re <= io_matrixIn_5_re; // @[R_Matrix_Estimation.scala 54:18]
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_x_reg_5_im <= 64'sh0; // @[R_Matrix_Estimation.scala 45:26]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      matrix_x_reg_5_im <= io_matrixIn_5_im; // @[R_Matrix_Estimation.scala 54:18]
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_x_reg_6_re <= 64'sh0; // @[R_Matrix_Estimation.scala 44:26]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      matrix_x_reg_6_re <= io_matrixIn_6_re; // @[R_Matrix_Estimation.scala 54:18]
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_x_reg_6_im <= 64'sh0; // @[R_Matrix_Estimation.scala 45:26]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      matrix_x_reg_6_im <= io_matrixIn_6_im; // @[R_Matrix_Estimation.scala 54:18]
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_x_reg_7_re <= 64'sh0; // @[R_Matrix_Estimation.scala 44:26]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      matrix_x_reg_7_re <= io_matrixIn_7_re; // @[R_Matrix_Estimation.scala 54:18]
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_x_reg_7_im <= 64'sh0; // @[R_Matrix_Estimation.scala 45:26]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      matrix_x_reg_7_im <= io_matrixIn_7_im; // @[R_Matrix_Estimation.scala 54:18]
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_0_re <= 64'sh0; // @[R_Matrix_Estimation.scala 48:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_0_re <= _GEN_131;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_0_im <= 64'sh0; // @[R_Matrix_Estimation.scala 49:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_0_im <= _GEN_130;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_1_re <= 64'sh0; // @[R_Matrix_Estimation.scala 48:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_1_re <= _GEN_133;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_1_im <= 64'sh0; // @[R_Matrix_Estimation.scala 49:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_1_im <= _GEN_132;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_2_re <= 64'sh0; // @[R_Matrix_Estimation.scala 48:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_2_re <= _GEN_135;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_2_im <= 64'sh0; // @[R_Matrix_Estimation.scala 49:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_2_im <= _GEN_134;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_3_re <= 64'sh0; // @[R_Matrix_Estimation.scala 48:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_3_re <= _GEN_137;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_3_im <= 64'sh0; // @[R_Matrix_Estimation.scala 49:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_3_im <= _GEN_136;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_4_re <= 64'sh0; // @[R_Matrix_Estimation.scala 48:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_4_re <= _GEN_139;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_4_im <= 64'sh0; // @[R_Matrix_Estimation.scala 49:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_4_im <= _GEN_138;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_5_re <= 64'sh0; // @[R_Matrix_Estimation.scala 48:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_5_re <= _GEN_141;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_5_im <= 64'sh0; // @[R_Matrix_Estimation.scala 49:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_5_im <= _GEN_140;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_6_re <= 64'sh0; // @[R_Matrix_Estimation.scala 48:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_6_re <= _GEN_143;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_6_im <= 64'sh0; // @[R_Matrix_Estimation.scala 49:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_6_im <= _GEN_142;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_7_re <= 64'sh0; // @[R_Matrix_Estimation.scala 48:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_7_re <= _GEN_145;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_7_im <= 64'sh0; // @[R_Matrix_Estimation.scala 49:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_7_im <= _GEN_144;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_8_re <= 64'sh0; // @[R_Matrix_Estimation.scala 48:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_8_re <= _GEN_147;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_8_im <= 64'sh0; // @[R_Matrix_Estimation.scala 49:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_8_im <= _GEN_146;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_9_re <= 64'sh0; // @[R_Matrix_Estimation.scala 48:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_9_re <= _GEN_149;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_9_im <= 64'sh0; // @[R_Matrix_Estimation.scala 49:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_9_im <= _GEN_148;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_10_re <= 64'sh0; // @[R_Matrix_Estimation.scala 48:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_10_re <= _GEN_151;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_10_im <= 64'sh0; // @[R_Matrix_Estimation.scala 49:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_10_im <= _GEN_150;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_11_re <= 64'sh0; // @[R_Matrix_Estimation.scala 48:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_11_re <= _GEN_153;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_11_im <= 64'sh0; // @[R_Matrix_Estimation.scala 49:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_11_im <= _GEN_152;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_12_re <= 64'sh0; // @[R_Matrix_Estimation.scala 48:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_12_re <= _GEN_155;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_12_im <= 64'sh0; // @[R_Matrix_Estimation.scala 49:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_12_im <= _GEN_154;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_13_re <= 64'sh0; // @[R_Matrix_Estimation.scala 48:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_13_re <= _GEN_157;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_13_im <= 64'sh0; // @[R_Matrix_Estimation.scala 49:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_13_im <= _GEN_156;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_14_re <= 64'sh0; // @[R_Matrix_Estimation.scala 48:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_14_re <= _GEN_159;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_14_im <= 64'sh0; // @[R_Matrix_Estimation.scala 49:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_14_im <= _GEN_158;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_15_re <= 64'sh0; // @[R_Matrix_Estimation.scala 48:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_15_re <= _GEN_161;
        end
      end
    end
    if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      matrix_mul_res_reg_15_im <= 64'sh0; // @[R_Matrix_Estimation.scala 49:32]
    end else if (!(io_ready)) begin // @[R_Matrix_Estimation.scala 53:24]
      if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
        if (status == 8'h2) begin // @[R_Matrix_Estimation.scala 67:32]
          matrix_mul_res_reg_15_im <= _GEN_160;
        end
      end
    end
    if (reset) begin // @[R_Matrix_Estimation.scala 30:29]
      status <= 8'h0; // @[R_Matrix_Estimation.scala 30:29]
    end else if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      status <= 8'h0; // @[R_Matrix_Estimation.scala 51:12]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      status <= 8'h1; // @[R_Matrix_Estimation.scala 55:12]
    end else if (status == 8'h1) begin // @[R_Matrix_Estimation.scala 58:26]
      status <= 8'h2; // @[R_Matrix_Estimation.scala 66:14]
    end else begin
      status <= _GEN_232;
    end
    if (reset) begin // @[R_Matrix_Estimation.scala 31:30]
      mul_cnt <= 3'h0; // @[R_Matrix_Estimation.scala 31:30]
    end else if (io_reset) begin // @[R_Matrix_Estimation.scala 42:18]
      mul_cnt <= 3'h0; // @[R_Matrix_Estimation.scala 52:13]
    end else if (io_ready) begin // @[R_Matrix_Estimation.scala 53:24]
      mul_cnt <= 3'h0; // @[R_Matrix_Estimation.scala 56:13]
    end else if (!(status == 8'h1)) begin // @[R_Matrix_Estimation.scala 58:26]
      mul_cnt <= _GEN_233;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  matrix_x_reg_0_re = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  matrix_x_reg_0_im = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  matrix_x_reg_1_re = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  matrix_x_reg_1_im = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  matrix_x_reg_2_re = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  matrix_x_reg_2_im = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  matrix_x_reg_3_re = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  matrix_x_reg_3_im = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  matrix_x_reg_4_re = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  matrix_x_reg_4_im = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  matrix_x_reg_5_re = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  matrix_x_reg_5_im = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  matrix_x_reg_6_re = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  matrix_x_reg_6_im = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  matrix_x_reg_7_re = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  matrix_x_reg_7_im = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  matrix_mul_res_reg_0_re = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  matrix_mul_res_reg_0_im = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  matrix_mul_res_reg_1_re = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  matrix_mul_res_reg_1_im = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  matrix_mul_res_reg_2_re = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  matrix_mul_res_reg_2_im = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  matrix_mul_res_reg_3_re = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  matrix_mul_res_reg_3_im = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  matrix_mul_res_reg_4_re = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  matrix_mul_res_reg_4_im = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  matrix_mul_res_reg_5_re = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  matrix_mul_res_reg_5_im = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  matrix_mul_res_reg_6_re = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  matrix_mul_res_reg_6_im = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  matrix_mul_res_reg_7_re = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  matrix_mul_res_reg_7_im = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  matrix_mul_res_reg_8_re = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  matrix_mul_res_reg_8_im = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  matrix_mul_res_reg_9_re = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  matrix_mul_res_reg_9_im = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  matrix_mul_res_reg_10_re = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  matrix_mul_res_reg_10_im = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  matrix_mul_res_reg_11_re = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  matrix_mul_res_reg_11_im = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  matrix_mul_res_reg_12_re = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  matrix_mul_res_reg_12_im = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  matrix_mul_res_reg_13_re = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  matrix_mul_res_reg_13_im = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  matrix_mul_res_reg_14_re = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  matrix_mul_res_reg_14_im = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  matrix_mul_res_reg_15_re = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  matrix_mul_res_reg_15_im = _RAND_47[63:0];
  _RAND_48 = {1{`RANDOM}};
  status = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  mul_cnt = _RAND_49[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module shift_range_1_8(
  input  [63:0] io_x,
  output [63:0] io_out,
  output [7:0]  io_cnt
);
  wire  _T = $signed(io_x) < 64'sh100000000; // @[Cordic_HV_Square_Root.scala 80:15]
  wire  index__0 = _T ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 84:90 85:18 87:18]
  wire [65:0] _T_3 = {$signed(io_x), 2'h0}; // @[Cordic_HV_Square_Root.scala 84:20]
  wire  index__1 = $signed(_T_3) < 66'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 84:90 85:18 87:18]
  wire [67:0] _T_5 = {$signed(io_x), 4'h0}; // @[Cordic_HV_Square_Root.scala 84:20]
  wire  index__2 = $signed(_T_5) < 68'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 84:90 85:18 87:18]
  wire [69:0] _T_7 = {$signed(io_x), 6'h0}; // @[Cordic_HV_Square_Root.scala 84:20]
  wire  index__3 = $signed(_T_7) < 70'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 84:90 85:18 87:18]
  wire [71:0] _T_9 = {$signed(io_x), 8'h0}; // @[Cordic_HV_Square_Root.scala 84:20]
  wire  index__4 = $signed(_T_9) < 72'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 84:90 85:18 87:18]
  wire [73:0] _T_11 = {$signed(io_x), 10'h0}; // @[Cordic_HV_Square_Root.scala 84:20]
  wire  index__5 = $signed(_T_11) < 74'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 84:90 85:18 87:18]
  wire [75:0] _T_13 = {$signed(io_x), 12'h0}; // @[Cordic_HV_Square_Root.scala 84:20]
  wire  index__6 = $signed(_T_13) < 76'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 84:90 85:18 87:18]
  wire [77:0] _T_15 = {$signed(io_x), 14'h0}; // @[Cordic_HV_Square_Root.scala 84:20]
  wire  index__7 = $signed(_T_15) < 78'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 84:90 85:18 87:18]
  wire [79:0] _T_17 = {$signed(io_x), 16'h0}; // @[Cordic_HV_Square_Root.scala 84:20]
  wire  index__8 = $signed(_T_17) < 80'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 84:90 85:18 87:18]
  wire [81:0] _T_19 = {$signed(io_x), 18'h0}; // @[Cordic_HV_Square_Root.scala 84:20]
  wire  index__9 = $signed(_T_19) < 82'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 84:90 85:18 87:18]
  wire [83:0] _T_21 = {$signed(io_x), 20'h0}; // @[Cordic_HV_Square_Root.scala 84:20]
  wire  index__10 = $signed(_T_21) < 84'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 84:90 85:18 87:18]
  wire [85:0] _T_23 = {$signed(io_x), 22'h0}; // @[Cordic_HV_Square_Root.scala 84:20]
  wire  index__11 = $signed(_T_23) < 86'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 84:90 85:18 87:18]
  wire [87:0] _T_25 = {$signed(io_x), 24'h0}; // @[Cordic_HV_Square_Root.scala 84:20]
  wire  index__12 = $signed(_T_25) < 88'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 84:90 85:18 87:18]
  wire [89:0] _T_27 = {$signed(io_x), 26'h0}; // @[Cordic_HV_Square_Root.scala 84:20]
  wire  index__13 = $signed(_T_27) < 90'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 84:90 85:18 87:18]
  wire [91:0] _T_29 = {$signed(io_x), 28'h0}; // @[Cordic_HV_Square_Root.scala 84:20]
  wire  index__14 = $signed(_T_29) < 92'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 84:90 85:18 87:18]
  wire [93:0] _T_31 = {$signed(io_x), 30'h0}; // @[Cordic_HV_Square_Root.scala 84:20]
  wire  index__15 = $signed(_T_31) < 94'sh100000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 84:90 85:18 87:18]
  wire [7:0] temp_cnt_lo = {index__7,index__6,index__5,index__4,index__3,index__2,index__1,index__0}; // @[Cordic_HV_Square_Root.scala 91:48]
  wire [15:0] _temp_cnt_T = {index__15,index__14,index__13,index__12,index__11,index__10,index__9,index__8,temp_cnt_lo}; // @[Cordic_HV_Square_Root.scala 91:48]
  wire [3:0] _temp_cnt_T_17 = _temp_cnt_T[14] ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_18 = _temp_cnt_T[13] ? 4'hd : _temp_cnt_T_17; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_19 = _temp_cnt_T[12] ? 4'hc : _temp_cnt_T_18; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_20 = _temp_cnt_T[11] ? 4'hb : _temp_cnt_T_19; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_21 = _temp_cnt_T[10] ? 4'ha : _temp_cnt_T_20; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_22 = _temp_cnt_T[9] ? 4'h9 : _temp_cnt_T_21; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_23 = _temp_cnt_T[8] ? 4'h8 : _temp_cnt_T_22; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_24 = _temp_cnt_T[7] ? 4'h7 : _temp_cnt_T_23; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_25 = _temp_cnt_T[6] ? 4'h6 : _temp_cnt_T_24; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_26 = _temp_cnt_T[5] ? 4'h5 : _temp_cnt_T_25; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_27 = _temp_cnt_T[4] ? 4'h4 : _temp_cnt_T_26; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_28 = _temp_cnt_T[3] ? 4'h3 : _temp_cnt_T_27; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_29 = _temp_cnt_T[2] ? 4'h2 : _temp_cnt_T_28; // @[Mux.scala 47:70]
  wire [3:0] _temp_cnt_T_30 = _temp_cnt_T[1] ? 4'h1 : _temp_cnt_T_29; // @[Mux.scala 47:70]
  wire [3:0] temp_cnt = _temp_cnt_T[0] ? 4'h0 : _temp_cnt_T_30; // @[Mux.scala 47:70]
  wire [4:0] _temp_uint_cnt_T = {temp_cnt, 1'h0}; // @[Cordic_HV_Square_Root.scala 92:32]
  wire  _T_33 = $signed(io_x) > 64'sh800000000; // @[Cordic_HV_Square_Root.scala 95:21]
  wire [37:0] _T_60 = io_x[63:26]; // @[Cordic_HV_Square_Root.scala 99:20]
  wire [63:0] _GEN_54 = {{26{_T_60[37]}},_T_60}; // @[Cordic_HV_Square_Root.scala 99:33]
  wire  index_1_13 = $signed(_GEN_54) > 64'sh800000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 100:18 102:18 99:90]
  wire [39:0] _T_58 = io_x[63:24]; // @[Cordic_HV_Square_Root.scala 99:20]
  wire [63:0] _GEN_55 = {{24{_T_58[39]}},_T_58}; // @[Cordic_HV_Square_Root.scala 99:33]
  wire  index_1_12 = $signed(_GEN_55) > 64'sh800000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 100:18 102:18 99:90]
  wire [41:0] _T_56 = io_x[63:22]; // @[Cordic_HV_Square_Root.scala 99:20]
  wire [63:0] _GEN_56 = {{22{_T_56[41]}},_T_56}; // @[Cordic_HV_Square_Root.scala 99:33]
  wire  index_1_11 = $signed(_GEN_56) > 64'sh800000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 100:18 102:18 99:90]
  wire [43:0] _T_54 = io_x[63:20]; // @[Cordic_HV_Square_Root.scala 99:20]
  wire [63:0] _GEN_57 = {{20{_T_54[43]}},_T_54}; // @[Cordic_HV_Square_Root.scala 99:33]
  wire  index_1_10 = $signed(_GEN_57) > 64'sh800000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 100:18 102:18 99:90]
  wire [45:0] _T_52 = io_x[63:18]; // @[Cordic_HV_Square_Root.scala 99:20]
  wire [63:0] _GEN_58 = {{18{_T_52[45]}},_T_52}; // @[Cordic_HV_Square_Root.scala 99:33]
  wire  index_1_9 = $signed(_GEN_58) > 64'sh800000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 100:18 102:18 99:90]
  wire [47:0] _T_50 = io_x[63:16]; // @[Cordic_HV_Square_Root.scala 99:20]
  wire [63:0] _GEN_59 = {{16{_T_50[47]}},_T_50}; // @[Cordic_HV_Square_Root.scala 99:33]
  wire  index_1_8 = $signed(_GEN_59) > 64'sh800000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 100:18 102:18 99:90]
  wire [49:0] _T_48 = io_x[63:14]; // @[Cordic_HV_Square_Root.scala 99:20]
  wire [63:0] _GEN_60 = {{14{_T_48[49]}},_T_48}; // @[Cordic_HV_Square_Root.scala 99:33]
  wire  index_1_7 = $signed(_GEN_60) > 64'sh800000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 100:18 102:18 99:90]
  wire [51:0] _T_46 = io_x[63:12]; // @[Cordic_HV_Square_Root.scala 99:20]
  wire [63:0] _GEN_61 = {{12{_T_46[51]}},_T_46}; // @[Cordic_HV_Square_Root.scala 99:33]
  wire  index_1_6 = $signed(_GEN_61) > 64'sh800000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 100:18 102:18 99:90]
  wire [53:0] _T_44 = io_x[63:10]; // @[Cordic_HV_Square_Root.scala 99:20]
  wire [63:0] _GEN_62 = {{10{_T_44[53]}},_T_44}; // @[Cordic_HV_Square_Root.scala 99:33]
  wire  index_1_5 = $signed(_GEN_62) > 64'sh800000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 100:18 102:18 99:90]
  wire [55:0] _T_42 = io_x[63:8]; // @[Cordic_HV_Square_Root.scala 99:20]
  wire [63:0] _GEN_63 = {{8{_T_42[55]}},_T_42}; // @[Cordic_HV_Square_Root.scala 99:33]
  wire  index_1_4 = $signed(_GEN_63) > 64'sh800000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 100:18 102:18 99:90]
  wire [57:0] _T_40 = io_x[63:6]; // @[Cordic_HV_Square_Root.scala 99:20]
  wire [63:0] _GEN_64 = {{6{_T_40[57]}},_T_40}; // @[Cordic_HV_Square_Root.scala 99:33]
  wire  index_1_3 = $signed(_GEN_64) > 64'sh800000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 100:18 102:18 99:90]
  wire [59:0] _T_38 = io_x[63:4]; // @[Cordic_HV_Square_Root.scala 99:20]
  wire [63:0] _GEN_65 = {{4{_T_38[59]}},_T_38}; // @[Cordic_HV_Square_Root.scala 99:33]
  wire  index_1_2 = $signed(_GEN_65) > 64'sh800000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 100:18 102:18 99:90]
  wire [61:0] _T_36 = io_x[63:2]; // @[Cordic_HV_Square_Root.scala 99:20]
  wire [63:0] _GEN_66 = {{2{_T_36[61]}},_T_36}; // @[Cordic_HV_Square_Root.scala 99:33]
  wire  index_1_1 = $signed(_GEN_66) > 64'sh800000000 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 100:18 102:18 99:90]
  wire  index_1_0 = _T_33 ? 1'h0 : 1'h1; // @[Cordic_HV_Square_Root.scala 100:18 102:18 99:90]
  wire [7:0] temp_cnt_lo_lo_1 = {index_1_7,index_1_6,index_1_5,index_1_4,index_1_3,index_1_2,index_1_1,index_1_0}; // @[Cordic_HV_Square_Root.scala 106:48]
  wire [31:0] _temp_cnt_T_31 = {16'hffff,2'h3,index_1_13,index_1_12,index_1_11,index_1_10,index_1_9,index_1_8,
    temp_cnt_lo_lo_1}; // @[Cordic_HV_Square_Root.scala 106:48]
  wire [4:0] _temp_cnt_T_64 = _temp_cnt_T_31[30] ? 5'h1e : 5'h1f; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_65 = _temp_cnt_T_31[29] ? 5'h1d : _temp_cnt_T_64; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_66 = _temp_cnt_T_31[28] ? 5'h1c : _temp_cnt_T_65; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_67 = _temp_cnt_T_31[27] ? 5'h1b : _temp_cnt_T_66; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_68 = _temp_cnt_T_31[26] ? 5'h1a : _temp_cnt_T_67; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_69 = _temp_cnt_T_31[25] ? 5'h19 : _temp_cnt_T_68; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_70 = _temp_cnt_T_31[24] ? 5'h18 : _temp_cnt_T_69; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_71 = _temp_cnt_T_31[23] ? 5'h17 : _temp_cnt_T_70; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_72 = _temp_cnt_T_31[22] ? 5'h16 : _temp_cnt_T_71; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_73 = _temp_cnt_T_31[21] ? 5'h15 : _temp_cnt_T_72; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_74 = _temp_cnt_T_31[20] ? 5'h14 : _temp_cnt_T_73; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_75 = _temp_cnt_T_31[19] ? 5'h13 : _temp_cnt_T_74; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_76 = _temp_cnt_T_31[18] ? 5'h12 : _temp_cnt_T_75; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_77 = _temp_cnt_T_31[17] ? 5'h11 : _temp_cnt_T_76; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_78 = _temp_cnt_T_31[16] ? 5'h10 : _temp_cnt_T_77; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_79 = _temp_cnt_T_31[15] ? 5'hf : _temp_cnt_T_78; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_80 = _temp_cnt_T_31[14] ? 5'he : _temp_cnt_T_79; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_81 = _temp_cnt_T_31[13] ? 5'hd : _temp_cnt_T_80; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_82 = _temp_cnt_T_31[12] ? 5'hc : _temp_cnt_T_81; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_83 = _temp_cnt_T_31[11] ? 5'hb : _temp_cnt_T_82; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_84 = _temp_cnt_T_31[10] ? 5'ha : _temp_cnt_T_83; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_85 = _temp_cnt_T_31[9] ? 5'h9 : _temp_cnt_T_84; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_86 = _temp_cnt_T_31[8] ? 5'h8 : _temp_cnt_T_85; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_87 = _temp_cnt_T_31[7] ? 5'h7 : _temp_cnt_T_86; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_88 = _temp_cnt_T_31[6] ? 5'h6 : _temp_cnt_T_87; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_89 = _temp_cnt_T_31[5] ? 5'h5 : _temp_cnt_T_88; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_90 = _temp_cnt_T_31[4] ? 5'h4 : _temp_cnt_T_89; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_91 = _temp_cnt_T_31[3] ? 5'h3 : _temp_cnt_T_90; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_92 = _temp_cnt_T_31[2] ? 5'h2 : _temp_cnt_T_91; // @[Mux.scala 47:70]
  wire [4:0] _temp_cnt_T_93 = _temp_cnt_T_31[1] ? 5'h1 : _temp_cnt_T_92; // @[Mux.scala 47:70]
  wire [4:0] temp_cnt_1 = _temp_cnt_T_31[0] ? 5'h0 : _temp_cnt_T_93; // @[Mux.scala 47:70]
  wire [5:0] _temp_uint_cnt_T_1 = {temp_cnt_1, 1'h0}; // @[Cordic_HV_Square_Root.scala 107:32]
  wire [7:0] _GEN_48 = $signed(io_x) > 64'sh800000000 ? {{2'd0}, _temp_uint_cnt_T_1} : 8'h0; // @[Cordic_HV_Square_Root.scala 107:19 95:78]
  wire [7:0] _io_cnt_T = $signed(io_x) < 64'sh100000000 ? {{3'd0}, _temp_uint_cnt_T} : _GEN_48; // @[Cordic_HV_Square_Root.scala 93:35]
  wire [94:0] _GEN_0 = {{31{io_x[63]}},io_x}; // @[Cordic_HV_Square_Root.scala 94:25]
  wire [94:0] _temp_out_T_1 = $signed(_GEN_0) << _temp_uint_cnt_T; // @[Cordic_HV_Square_Root.scala 94:25]
  wire [7:0] _io_cnt_T_4 = 8'sh0 - $signed(_io_cnt_T); // @[Cordic_HV_Square_Root.scala 108:15]
  wire [63:0] _temp_out_T_3 = $signed(io_x) >>> _temp_uint_cnt_T_1; // @[Cordic_HV_Square_Root.scala 109:25]
  wire [7:0] _GEN_49 = $signed(io_x) > 64'sh800000000 ? $signed(_io_cnt_T_4) : $signed(8'sh0); // @[Cordic_HV_Square_Root.scala 108:12 111:12 95:78]
  wire [63:0] _GEN_50 = $signed(io_x) > 64'sh800000000 ? $signed(_temp_out_T_3) : $signed(io_x); // @[Cordic_HV_Square_Root.scala 109:14 112:14 95:78]
  wire [94:0] _GEN_53 = $signed(io_x) < 64'sh100000000 ? $signed(_temp_out_T_1) : $signed({{31{_GEN_50[63]}},_GEN_50}); // @[Cordic_HV_Square_Root.scala 80:72 94:14]
  assign io_out = _GEN_53[63:0]; // @[Cordic_HV_Square_Root.scala 77:34]
  assign io_cnt = $signed(io_x) < 64'sh100000000 ? $signed(_io_cnt_T) : $signed(_GEN_49); // @[Cordic_HV_Square_Root.scala 80:72 93:12]
endmodule
module cordic_hv_square_root_origin(
  input         clock,
  input         reset,
  input  [63:0] io_in,
  output [63:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] x = $signed(io_in) + 64'sh100000000; // @[Cordic_HV_Square_Root.scala 23:29]
  wire [63:0] y = $signed(io_in) - 64'sh100000000; // @[Cordic_HV_Square_Root.scala 24:29]
  reg [63:0] current_x_0; // @[Cordic_HV_Square_Root.scala 30:43]
  reg [63:0] current_x_1; // @[Cordic_HV_Square_Root.scala 30:43]
  reg [63:0] current_x_2; // @[Cordic_HV_Square_Root.scala 30:43]
  reg [63:0] current_x_3; // @[Cordic_HV_Square_Root.scala 30:43]
  reg [63:0] current_x_4; // @[Cordic_HV_Square_Root.scala 30:43]
  reg [63:0] current_x_5; // @[Cordic_HV_Square_Root.scala 30:43]
  reg [63:0] current_x_6; // @[Cordic_HV_Square_Root.scala 30:43]
  reg [63:0] current_x_7; // @[Cordic_HV_Square_Root.scala 30:43]
  reg [63:0] current_x_8; // @[Cordic_HV_Square_Root.scala 30:43]
  reg [63:0] current_x_9; // @[Cordic_HV_Square_Root.scala 30:43]
  reg [63:0] current_x_10; // @[Cordic_HV_Square_Root.scala 30:43]
  reg [63:0] current_x_11; // @[Cordic_HV_Square_Root.scala 30:43]
  reg [63:0] current_x_12; // @[Cordic_HV_Square_Root.scala 30:43]
  reg [63:0] current_x_13; // @[Cordic_HV_Square_Root.scala 30:43]
  reg [63:0] current_x_14; // @[Cordic_HV_Square_Root.scala 30:43]
  reg [63:0] current_y_0; // @[Cordic_HV_Square_Root.scala 31:43]
  reg [63:0] current_y_1; // @[Cordic_HV_Square_Root.scala 31:43]
  reg [63:0] current_y_2; // @[Cordic_HV_Square_Root.scala 31:43]
  reg [63:0] current_y_3; // @[Cordic_HV_Square_Root.scala 31:43]
  reg [63:0] current_y_4; // @[Cordic_HV_Square_Root.scala 31:43]
  reg [63:0] current_y_5; // @[Cordic_HV_Square_Root.scala 31:43]
  reg [63:0] current_y_6; // @[Cordic_HV_Square_Root.scala 31:43]
  reg [63:0] current_y_7; // @[Cordic_HV_Square_Root.scala 31:43]
  reg [63:0] current_y_8; // @[Cordic_HV_Square_Root.scala 31:43]
  reg [63:0] current_y_9; // @[Cordic_HV_Square_Root.scala 31:43]
  reg [63:0] current_y_10; // @[Cordic_HV_Square_Root.scala 31:43]
  reg [63:0] current_y_11; // @[Cordic_HV_Square_Root.scala 31:43]
  reg [63:0] current_y_12; // @[Cordic_HV_Square_Root.scala 31:43]
  reg [63:0] current_y_13; // @[Cordic_HV_Square_Root.scala 31:43]
  wire [62:0] _current_x_0_T = y[63:1]; // @[Cordic_HV_Square_Root.scala 42:36]
  wire [63:0] _GEN_30 = {{1{_current_x_0_T[62]}},_current_x_0_T}; // @[Cordic_HV_Square_Root.scala 42:31]
  wire [63:0] _current_x_0_T_3 = $signed(x) + $signed(_GEN_30); // @[Cordic_HV_Square_Root.scala 42:31]
  wire [62:0] _current_y_0_T = x[63:1]; // @[Cordic_HV_Square_Root.scala 43:36]
  wire [63:0] _GEN_31 = {{1{_current_y_0_T[62]}},_current_y_0_T}; // @[Cordic_HV_Square_Root.scala 43:31]
  wire [63:0] _current_y_0_T_3 = $signed(y) + $signed(_GEN_31); // @[Cordic_HV_Square_Root.scala 43:31]
  wire [63:0] _current_x_0_T_7 = $signed(x) - $signed(_GEN_30); // @[Cordic_HV_Square_Root.scala 45:31]
  wire [63:0] _current_y_0_T_7 = $signed(y) - $signed(_GEN_31); // @[Cordic_HV_Square_Root.scala 46:31]
  wire [61:0] _current_x_1_T = current_y_0[63:2]; // @[Cordic_HV_Square_Root.scala 50:66]
  wire [63:0] _GEN_34 = {{2{_current_x_1_T[61]}},_current_x_1_T}; // @[Cordic_HV_Square_Root.scala 50:46]
  wire [63:0] _current_x_1_T_3 = $signed(current_x_0) + $signed(_GEN_34); // @[Cordic_HV_Square_Root.scala 50:46]
  wire [61:0] _current_y_1_T = current_x_0[63:2]; // @[Cordic_HV_Square_Root.scala 51:66]
  wire [63:0] _GEN_35 = {{2{_current_y_1_T[61]}},_current_y_1_T}; // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_y_1_T_3 = $signed(current_y_0) + $signed(_GEN_35); // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_x_1_T_7 = $signed(current_x_0) - $signed(_GEN_34); // @[Cordic_HV_Square_Root.scala 53:46]
  wire [63:0] _current_y_1_T_7 = $signed(current_y_0) - $signed(_GEN_35); // @[Cordic_HV_Square_Root.scala 54:46]
  wire [60:0] _current_x_2_T = current_y_1[63:3]; // @[Cordic_HV_Square_Root.scala 50:66]
  wire [63:0] _GEN_38 = {{3{_current_x_2_T[60]}},_current_x_2_T}; // @[Cordic_HV_Square_Root.scala 50:46]
  wire [63:0] _current_x_2_T_3 = $signed(current_x_1) + $signed(_GEN_38); // @[Cordic_HV_Square_Root.scala 50:46]
  wire [60:0] _current_y_2_T = current_x_1[63:3]; // @[Cordic_HV_Square_Root.scala 51:66]
  wire [63:0] _GEN_39 = {{3{_current_y_2_T[60]}},_current_y_2_T}; // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_y_2_T_3 = $signed(current_y_1) + $signed(_GEN_39); // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_x_2_T_7 = $signed(current_x_1) - $signed(_GEN_38); // @[Cordic_HV_Square_Root.scala 53:46]
  wire [63:0] _current_y_2_T_7 = $signed(current_y_1) - $signed(_GEN_39); // @[Cordic_HV_Square_Root.scala 54:46]
  wire [59:0] _current_x_3_T = current_y_2[63:4]; // @[Cordic_HV_Square_Root.scala 50:66]
  wire [63:0] _GEN_42 = {{4{_current_x_3_T[59]}},_current_x_3_T}; // @[Cordic_HV_Square_Root.scala 50:46]
  wire [63:0] _current_x_3_T_3 = $signed(current_x_2) + $signed(_GEN_42); // @[Cordic_HV_Square_Root.scala 50:46]
  wire [59:0] _current_y_3_T = current_x_2[63:4]; // @[Cordic_HV_Square_Root.scala 51:66]
  wire [63:0] _GEN_43 = {{4{_current_y_3_T[59]}},_current_y_3_T}; // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_y_3_T_3 = $signed(current_y_2) + $signed(_GEN_43); // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_x_3_T_7 = $signed(current_x_2) - $signed(_GEN_42); // @[Cordic_HV_Square_Root.scala 53:46]
  wire [63:0] _current_y_3_T_7 = $signed(current_y_2) - $signed(_GEN_43); // @[Cordic_HV_Square_Root.scala 54:46]
  wire [58:0] _current_x_4_T = current_y_3[63:5]; // @[Cordic_HV_Square_Root.scala 50:66]
  wire [63:0] _GEN_46 = {{5{_current_x_4_T[58]}},_current_x_4_T}; // @[Cordic_HV_Square_Root.scala 50:46]
  wire [63:0] _current_x_4_T_3 = $signed(current_x_3) + $signed(_GEN_46); // @[Cordic_HV_Square_Root.scala 50:46]
  wire [58:0] _current_y_4_T = current_x_3[63:5]; // @[Cordic_HV_Square_Root.scala 51:66]
  wire [63:0] _GEN_47 = {{5{_current_y_4_T[58]}},_current_y_4_T}; // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_y_4_T_3 = $signed(current_y_3) + $signed(_GEN_47); // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_x_4_T_7 = $signed(current_x_3) - $signed(_GEN_46); // @[Cordic_HV_Square_Root.scala 53:46]
  wire [63:0] _current_y_4_T_7 = $signed(current_y_3) - $signed(_GEN_47); // @[Cordic_HV_Square_Root.scala 54:46]
  wire [57:0] _current_x_5_T = current_y_4[63:6]; // @[Cordic_HV_Square_Root.scala 50:66]
  wire [63:0] _GEN_50 = {{6{_current_x_5_T[57]}},_current_x_5_T}; // @[Cordic_HV_Square_Root.scala 50:46]
  wire [63:0] _current_x_5_T_3 = $signed(current_x_4) + $signed(_GEN_50); // @[Cordic_HV_Square_Root.scala 50:46]
  wire [57:0] _current_y_5_T = current_x_4[63:6]; // @[Cordic_HV_Square_Root.scala 51:66]
  wire [63:0] _GEN_51 = {{6{_current_y_5_T[57]}},_current_y_5_T}; // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_y_5_T_3 = $signed(current_y_4) + $signed(_GEN_51); // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_x_5_T_7 = $signed(current_x_4) - $signed(_GEN_50); // @[Cordic_HV_Square_Root.scala 53:46]
  wire [63:0] _current_y_5_T_7 = $signed(current_y_4) - $signed(_GEN_51); // @[Cordic_HV_Square_Root.scala 54:46]
  wire [56:0] _current_x_6_T = current_y_5[63:7]; // @[Cordic_HV_Square_Root.scala 50:66]
  wire [63:0] _GEN_54 = {{7{_current_x_6_T[56]}},_current_x_6_T}; // @[Cordic_HV_Square_Root.scala 50:46]
  wire [63:0] _current_x_6_T_3 = $signed(current_x_5) + $signed(_GEN_54); // @[Cordic_HV_Square_Root.scala 50:46]
  wire [56:0] _current_y_6_T = current_x_5[63:7]; // @[Cordic_HV_Square_Root.scala 51:66]
  wire [63:0] _GEN_55 = {{7{_current_y_6_T[56]}},_current_y_6_T}; // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_y_6_T_3 = $signed(current_y_5) + $signed(_GEN_55); // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_x_6_T_7 = $signed(current_x_5) - $signed(_GEN_54); // @[Cordic_HV_Square_Root.scala 53:46]
  wire [63:0] _current_y_6_T_7 = $signed(current_y_5) - $signed(_GEN_55); // @[Cordic_HV_Square_Root.scala 54:46]
  wire [55:0] _current_x_7_T = current_y_6[63:8]; // @[Cordic_HV_Square_Root.scala 50:66]
  wire [63:0] _GEN_58 = {{8{_current_x_7_T[55]}},_current_x_7_T}; // @[Cordic_HV_Square_Root.scala 50:46]
  wire [63:0] _current_x_7_T_3 = $signed(current_x_6) + $signed(_GEN_58); // @[Cordic_HV_Square_Root.scala 50:46]
  wire [55:0] _current_y_7_T = current_x_6[63:8]; // @[Cordic_HV_Square_Root.scala 51:66]
  wire [63:0] _GEN_59 = {{8{_current_y_7_T[55]}},_current_y_7_T}; // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_y_7_T_3 = $signed(current_y_6) + $signed(_GEN_59); // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_x_7_T_7 = $signed(current_x_6) - $signed(_GEN_58); // @[Cordic_HV_Square_Root.scala 53:46]
  wire [63:0] _current_y_7_T_7 = $signed(current_y_6) - $signed(_GEN_59); // @[Cordic_HV_Square_Root.scala 54:46]
  wire [54:0] _current_x_8_T = current_y_7[63:9]; // @[Cordic_HV_Square_Root.scala 50:66]
  wire [63:0] _GEN_62 = {{9{_current_x_8_T[54]}},_current_x_8_T}; // @[Cordic_HV_Square_Root.scala 50:46]
  wire [63:0] _current_x_8_T_3 = $signed(current_x_7) + $signed(_GEN_62); // @[Cordic_HV_Square_Root.scala 50:46]
  wire [54:0] _current_y_8_T = current_x_7[63:9]; // @[Cordic_HV_Square_Root.scala 51:66]
  wire [63:0] _GEN_63 = {{9{_current_y_8_T[54]}},_current_y_8_T}; // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_y_8_T_3 = $signed(current_y_7) + $signed(_GEN_63); // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_x_8_T_7 = $signed(current_x_7) - $signed(_GEN_62); // @[Cordic_HV_Square_Root.scala 53:46]
  wire [63:0] _current_y_8_T_7 = $signed(current_y_7) - $signed(_GEN_63); // @[Cordic_HV_Square_Root.scala 54:46]
  wire [53:0] _current_x_9_T = current_y_8[63:10]; // @[Cordic_HV_Square_Root.scala 50:66]
  wire [63:0] _GEN_66 = {{10{_current_x_9_T[53]}},_current_x_9_T}; // @[Cordic_HV_Square_Root.scala 50:46]
  wire [63:0] _current_x_9_T_3 = $signed(current_x_8) + $signed(_GEN_66); // @[Cordic_HV_Square_Root.scala 50:46]
  wire [53:0] _current_y_9_T = current_x_8[63:10]; // @[Cordic_HV_Square_Root.scala 51:66]
  wire [63:0] _GEN_67 = {{10{_current_y_9_T[53]}},_current_y_9_T}; // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_y_9_T_3 = $signed(current_y_8) + $signed(_GEN_67); // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_x_9_T_7 = $signed(current_x_8) - $signed(_GEN_66); // @[Cordic_HV_Square_Root.scala 53:46]
  wire [63:0] _current_y_9_T_7 = $signed(current_y_8) - $signed(_GEN_67); // @[Cordic_HV_Square_Root.scala 54:46]
  wire [52:0] _current_x_10_T = current_y_9[63:11]; // @[Cordic_HV_Square_Root.scala 50:66]
  wire [63:0] _GEN_70 = {{11{_current_x_10_T[52]}},_current_x_10_T}; // @[Cordic_HV_Square_Root.scala 50:46]
  wire [63:0] _current_x_10_T_3 = $signed(current_x_9) + $signed(_GEN_70); // @[Cordic_HV_Square_Root.scala 50:46]
  wire [52:0] _current_y_10_T = current_x_9[63:11]; // @[Cordic_HV_Square_Root.scala 51:66]
  wire [63:0] _GEN_71 = {{11{_current_y_10_T[52]}},_current_y_10_T}; // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_y_10_T_3 = $signed(current_y_9) + $signed(_GEN_71); // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_x_10_T_7 = $signed(current_x_9) - $signed(_GEN_70); // @[Cordic_HV_Square_Root.scala 53:46]
  wire [63:0] _current_y_10_T_7 = $signed(current_y_9) - $signed(_GEN_71); // @[Cordic_HV_Square_Root.scala 54:46]
  wire [51:0] _current_x_11_T = current_y_10[63:12]; // @[Cordic_HV_Square_Root.scala 50:66]
  wire [63:0] _GEN_74 = {{12{_current_x_11_T[51]}},_current_x_11_T}; // @[Cordic_HV_Square_Root.scala 50:46]
  wire [63:0] _current_x_11_T_3 = $signed(current_x_10) + $signed(_GEN_74); // @[Cordic_HV_Square_Root.scala 50:46]
  wire [51:0] _current_y_11_T = current_x_10[63:12]; // @[Cordic_HV_Square_Root.scala 51:66]
  wire [63:0] _GEN_75 = {{12{_current_y_11_T[51]}},_current_y_11_T}; // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_y_11_T_3 = $signed(current_y_10) + $signed(_GEN_75); // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_x_11_T_7 = $signed(current_x_10) - $signed(_GEN_74); // @[Cordic_HV_Square_Root.scala 53:46]
  wire [63:0] _current_y_11_T_7 = $signed(current_y_10) - $signed(_GEN_75); // @[Cordic_HV_Square_Root.scala 54:46]
  wire [50:0] _current_x_12_T = current_y_11[63:13]; // @[Cordic_HV_Square_Root.scala 50:66]
  wire [63:0] _GEN_78 = {{13{_current_x_12_T[50]}},_current_x_12_T}; // @[Cordic_HV_Square_Root.scala 50:46]
  wire [63:0] _current_x_12_T_3 = $signed(current_x_11) + $signed(_GEN_78); // @[Cordic_HV_Square_Root.scala 50:46]
  wire [50:0] _current_y_12_T = current_x_11[63:13]; // @[Cordic_HV_Square_Root.scala 51:66]
  wire [63:0] _GEN_79 = {{13{_current_y_12_T[50]}},_current_y_12_T}; // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_y_12_T_3 = $signed(current_y_11) + $signed(_GEN_79); // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_x_12_T_7 = $signed(current_x_11) - $signed(_GEN_78); // @[Cordic_HV_Square_Root.scala 53:46]
  wire [63:0] _current_y_12_T_7 = $signed(current_y_11) - $signed(_GEN_79); // @[Cordic_HV_Square_Root.scala 54:46]
  wire [49:0] _current_x_13_T = current_y_12[63:14]; // @[Cordic_HV_Square_Root.scala 50:66]
  wire [63:0] _GEN_82 = {{14{_current_x_13_T[49]}},_current_x_13_T}; // @[Cordic_HV_Square_Root.scala 50:46]
  wire [63:0] _current_x_13_T_3 = $signed(current_x_12) + $signed(_GEN_82); // @[Cordic_HV_Square_Root.scala 50:46]
  wire [49:0] _current_y_13_T = current_x_12[63:14]; // @[Cordic_HV_Square_Root.scala 51:66]
  wire [63:0] _GEN_83 = {{14{_current_y_13_T[49]}},_current_y_13_T}; // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_y_13_T_3 = $signed(current_y_12) + $signed(_GEN_83); // @[Cordic_HV_Square_Root.scala 51:46]
  wire [63:0] _current_x_13_T_7 = $signed(current_x_12) - $signed(_GEN_82); // @[Cordic_HV_Square_Root.scala 53:46]
  wire [63:0] _current_y_13_T_7 = $signed(current_y_12) - $signed(_GEN_83); // @[Cordic_HV_Square_Root.scala 54:46]
  wire [48:0] _current_x_14_T = current_y_13[63:15]; // @[Cordic_HV_Square_Root.scala 50:66]
  wire [63:0] _GEN_86 = {{15{_current_x_14_T[48]}},_current_x_14_T}; // @[Cordic_HV_Square_Root.scala 50:46]
  wire [63:0] _current_x_14_T_3 = $signed(current_x_13) + $signed(_GEN_86); // @[Cordic_HV_Square_Root.scala 50:46]
  wire [63:0] _current_x_14_T_7 = $signed(current_x_13) - $signed(_GEN_86); // @[Cordic_HV_Square_Root.scala 53:46]
  wire [127:0] _io_out_T = $signed(current_x_14) * 64'sh13483d0ff; // @[Cordic_HV_Square_Root.scala 59:44]
  wire [126:0] _io_out_T_1 = _io_out_T[127:1]; // @[Cordic_HV_Square_Root.scala 59:58]
  wire [94:0] _GEN_90 = _io_out_T_1[126:32]; // @[Cordic_HV_Square_Root.scala 59:10]
  assign io_out = _GEN_90[63:0]; // @[Cordic_HV_Square_Root.scala 59:10]
  always @(posedge clock) begin
    if (reset) begin // @[Cordic_HV_Square_Root.scala 30:43]
      current_x_0 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 30:43]
    end else if ($signed(y) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 41:73]
      current_x_0 <= _current_x_0_T_3; // @[Cordic_HV_Square_Root.scala 42:26]
    end else begin
      current_x_0 <= _current_x_0_T_7; // @[Cordic_HV_Square_Root.scala 45:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 30:43]
      current_x_1 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 30:43]
    end else if ($signed(current_y_0) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_x_1 <= _current_x_1_T_3; // @[Cordic_HV_Square_Root.scala 50:26]
    end else begin
      current_x_1 <= _current_x_1_T_7; // @[Cordic_HV_Square_Root.scala 53:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 30:43]
      current_x_2 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 30:43]
    end else if ($signed(current_y_1) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_x_2 <= _current_x_2_T_3; // @[Cordic_HV_Square_Root.scala 50:26]
    end else begin
      current_x_2 <= _current_x_2_T_7; // @[Cordic_HV_Square_Root.scala 53:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 30:43]
      current_x_3 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 30:43]
    end else if ($signed(current_y_2) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_x_3 <= _current_x_3_T_3; // @[Cordic_HV_Square_Root.scala 50:26]
    end else begin
      current_x_3 <= _current_x_3_T_7; // @[Cordic_HV_Square_Root.scala 53:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 30:43]
      current_x_4 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 30:43]
    end else if ($signed(current_y_3) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_x_4 <= _current_x_4_T_3; // @[Cordic_HV_Square_Root.scala 50:26]
    end else begin
      current_x_4 <= _current_x_4_T_7; // @[Cordic_HV_Square_Root.scala 53:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 30:43]
      current_x_5 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 30:43]
    end else if ($signed(current_y_4) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_x_5 <= _current_x_5_T_3; // @[Cordic_HV_Square_Root.scala 50:26]
    end else begin
      current_x_5 <= _current_x_5_T_7; // @[Cordic_HV_Square_Root.scala 53:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 30:43]
      current_x_6 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 30:43]
    end else if ($signed(current_y_5) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_x_6 <= _current_x_6_T_3; // @[Cordic_HV_Square_Root.scala 50:26]
    end else begin
      current_x_6 <= _current_x_6_T_7; // @[Cordic_HV_Square_Root.scala 53:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 30:43]
      current_x_7 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 30:43]
    end else if ($signed(current_y_6) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_x_7 <= _current_x_7_T_3; // @[Cordic_HV_Square_Root.scala 50:26]
    end else begin
      current_x_7 <= _current_x_7_T_7; // @[Cordic_HV_Square_Root.scala 53:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 30:43]
      current_x_8 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 30:43]
    end else if ($signed(current_y_7) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_x_8 <= _current_x_8_T_3; // @[Cordic_HV_Square_Root.scala 50:26]
    end else begin
      current_x_8 <= _current_x_8_T_7; // @[Cordic_HV_Square_Root.scala 53:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 30:43]
      current_x_9 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 30:43]
    end else if ($signed(current_y_8) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_x_9 <= _current_x_9_T_3; // @[Cordic_HV_Square_Root.scala 50:26]
    end else begin
      current_x_9 <= _current_x_9_T_7; // @[Cordic_HV_Square_Root.scala 53:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 30:43]
      current_x_10 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 30:43]
    end else if ($signed(current_y_9) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_x_10 <= _current_x_10_T_3; // @[Cordic_HV_Square_Root.scala 50:26]
    end else begin
      current_x_10 <= _current_x_10_T_7; // @[Cordic_HV_Square_Root.scala 53:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 30:43]
      current_x_11 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 30:43]
    end else if ($signed(current_y_10) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_x_11 <= _current_x_11_T_3; // @[Cordic_HV_Square_Root.scala 50:26]
    end else begin
      current_x_11 <= _current_x_11_T_7; // @[Cordic_HV_Square_Root.scala 53:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 30:43]
      current_x_12 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 30:43]
    end else if ($signed(current_y_11) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_x_12 <= _current_x_12_T_3; // @[Cordic_HV_Square_Root.scala 50:26]
    end else begin
      current_x_12 <= _current_x_12_T_7; // @[Cordic_HV_Square_Root.scala 53:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 30:43]
      current_x_13 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 30:43]
    end else if ($signed(current_y_12) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_x_13 <= _current_x_13_T_3; // @[Cordic_HV_Square_Root.scala 50:26]
    end else begin
      current_x_13 <= _current_x_13_T_7; // @[Cordic_HV_Square_Root.scala 53:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 30:43]
      current_x_14 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 30:43]
    end else if ($signed(current_y_13) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_x_14 <= _current_x_14_T_3; // @[Cordic_HV_Square_Root.scala 50:26]
    end else begin
      current_x_14 <= _current_x_14_T_7; // @[Cordic_HV_Square_Root.scala 53:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 31:43]
      current_y_0 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 31:43]
    end else if ($signed(y) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 41:73]
      current_y_0 <= _current_y_0_T_3; // @[Cordic_HV_Square_Root.scala 43:26]
    end else begin
      current_y_0 <= _current_y_0_T_7; // @[Cordic_HV_Square_Root.scala 46:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 31:43]
      current_y_1 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 31:43]
    end else if ($signed(current_y_0) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_y_1 <= _current_y_1_T_3; // @[Cordic_HV_Square_Root.scala 51:26]
    end else begin
      current_y_1 <= _current_y_1_T_7; // @[Cordic_HV_Square_Root.scala 54:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 31:43]
      current_y_2 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 31:43]
    end else if ($signed(current_y_1) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_y_2 <= _current_y_2_T_3; // @[Cordic_HV_Square_Root.scala 51:26]
    end else begin
      current_y_2 <= _current_y_2_T_7; // @[Cordic_HV_Square_Root.scala 54:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 31:43]
      current_y_3 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 31:43]
    end else if ($signed(current_y_2) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_y_3 <= _current_y_3_T_3; // @[Cordic_HV_Square_Root.scala 51:26]
    end else begin
      current_y_3 <= _current_y_3_T_7; // @[Cordic_HV_Square_Root.scala 54:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 31:43]
      current_y_4 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 31:43]
    end else if ($signed(current_y_3) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_y_4 <= _current_y_4_T_3; // @[Cordic_HV_Square_Root.scala 51:26]
    end else begin
      current_y_4 <= _current_y_4_T_7; // @[Cordic_HV_Square_Root.scala 54:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 31:43]
      current_y_5 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 31:43]
    end else if ($signed(current_y_4) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_y_5 <= _current_y_5_T_3; // @[Cordic_HV_Square_Root.scala 51:26]
    end else begin
      current_y_5 <= _current_y_5_T_7; // @[Cordic_HV_Square_Root.scala 54:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 31:43]
      current_y_6 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 31:43]
    end else if ($signed(current_y_5) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_y_6 <= _current_y_6_T_3; // @[Cordic_HV_Square_Root.scala 51:26]
    end else begin
      current_y_6 <= _current_y_6_T_7; // @[Cordic_HV_Square_Root.scala 54:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 31:43]
      current_y_7 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 31:43]
    end else if ($signed(current_y_6) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_y_7 <= _current_y_7_T_3; // @[Cordic_HV_Square_Root.scala 51:26]
    end else begin
      current_y_7 <= _current_y_7_T_7; // @[Cordic_HV_Square_Root.scala 54:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 31:43]
      current_y_8 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 31:43]
    end else if ($signed(current_y_7) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_y_8 <= _current_y_8_T_3; // @[Cordic_HV_Square_Root.scala 51:26]
    end else begin
      current_y_8 <= _current_y_8_T_7; // @[Cordic_HV_Square_Root.scala 54:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 31:43]
      current_y_9 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 31:43]
    end else if ($signed(current_y_8) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_y_9 <= _current_y_9_T_3; // @[Cordic_HV_Square_Root.scala 51:26]
    end else begin
      current_y_9 <= _current_y_9_T_7; // @[Cordic_HV_Square_Root.scala 54:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 31:43]
      current_y_10 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 31:43]
    end else if ($signed(current_y_9) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_y_10 <= _current_y_10_T_3; // @[Cordic_HV_Square_Root.scala 51:26]
    end else begin
      current_y_10 <= _current_y_10_T_7; // @[Cordic_HV_Square_Root.scala 54:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 31:43]
      current_y_11 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 31:43]
    end else if ($signed(current_y_10) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_y_11 <= _current_y_11_T_3; // @[Cordic_HV_Square_Root.scala 51:26]
    end else begin
      current_y_11 <= _current_y_11_T_7; // @[Cordic_HV_Square_Root.scala 54:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 31:43]
      current_y_12 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 31:43]
    end else if ($signed(current_y_11) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_y_12 <= _current_y_12_T_3; // @[Cordic_HV_Square_Root.scala 51:26]
    end else begin
      current_y_12 <= _current_y_12_T_7; // @[Cordic_HV_Square_Root.scala 54:26]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 31:43]
      current_y_13 <= 64'sh0; // @[Cordic_HV_Square_Root.scala 31:43]
    end else if ($signed(current_y_12) < 64'sh0) begin // @[Cordic_HV_Square_Root.scala 49:88]
      current_y_13 <= _current_y_13_T_3; // @[Cordic_HV_Square_Root.scala 51:26]
    end else begin
      current_y_13 <= _current_y_13_T_7; // @[Cordic_HV_Square_Root.scala 54:26]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  current_x_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  current_x_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  current_x_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  current_x_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  current_x_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  current_x_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  current_x_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  current_x_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  current_x_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  current_x_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  current_x_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  current_x_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  current_x_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  current_x_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  current_x_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  current_y_0 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  current_y_1 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  current_y_2 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  current_y_3 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  current_y_4 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  current_y_5 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  current_y_6 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  current_y_7 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  current_y_8 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  current_y_9 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  current_y_10 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  current_y_11 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  current_y_12 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  current_y_13 = _RAND_28[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cordic_hv_square_root(
  input         clock,
  input         reset,
  input  [63:0] io_in,
  output [63:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] unit_io_x; // @[Cordic_HV_Square_Root.scala 130:22]
  wire [63:0] unit_io_out; // @[Cordic_HV_Square_Root.scala 130:22]
  wire [7:0] unit_io_cnt; // @[Cordic_HV_Square_Root.scala 130:22]
  wire  unit_1_clock; // @[Cordic_HV_Square_Root.scala 176:20]
  wire  unit_1_reset; // @[Cordic_HV_Square_Root.scala 176:20]
  wire [63:0] unit_1_io_in; // @[Cordic_HV_Square_Root.scala 176:20]
  wire [63:0] unit_1_io_out; // @[Cordic_HV_Square_Root.scala 176:20]
  wire  flag = $signed(io_in) >= 64'sh0; // @[Cordic_HV_Square_Root.scala 156:14]
  wire [63:0] _temp_in_T_2 = 64'sh0 - $signed(io_in); // @[Cordic_HV_Square_Root.scala 160:16]
  reg [7:0] cnt_reg_0; // @[Cordic_HV_Square_Root.scala 167:35]
  reg [7:0] cnt_reg_1; // @[Cordic_HV_Square_Root.scala 167:35]
  reg [7:0] cnt_reg_2; // @[Cordic_HV_Square_Root.scala 167:35]
  reg [7:0] cnt_reg_3; // @[Cordic_HV_Square_Root.scala 167:35]
  reg [7:0] cnt_reg_4; // @[Cordic_HV_Square_Root.scala 167:35]
  reg [7:0] cnt_reg_5; // @[Cordic_HV_Square_Root.scala 167:35]
  reg [7:0] cnt_reg_6; // @[Cordic_HV_Square_Root.scala 167:35]
  reg [7:0] cnt_reg_7; // @[Cordic_HV_Square_Root.scala 167:35]
  reg [7:0] cnt_reg_8; // @[Cordic_HV_Square_Root.scala 167:35]
  reg [7:0] cnt_reg_9; // @[Cordic_HV_Square_Root.scala 167:35]
  reg [7:0] cnt_reg_10; // @[Cordic_HV_Square_Root.scala 167:35]
  reg [7:0] cnt_reg_11; // @[Cordic_HV_Square_Root.scala 167:35]
  reg [7:0] cnt_reg_12; // @[Cordic_HV_Square_Root.scala 167:35]
  reg [7:0] cnt_reg_13; // @[Cordic_HV_Square_Root.scala 167:35]
  reg [7:0] cnt_reg_14; // @[Cordic_HV_Square_Root.scala 167:35]
  wire [7:0] u_cnt = cnt_reg_14; // @[Cordic_HV_Square_Root.scala 181:51]
  wire [63:0] _temp_out_T_1 = $signed(unit_1_io_out) >>> u_cnt[7:1]; // @[Cordic_HV_Square_Root.scala 182:30]
  wire [7:0] u_cnt_1 = 8'sh0 - $signed(cnt_reg_14); // @[Cordic_HV_Square_Root.scala 184:54]
  wire [190:0] _GEN_0 = {{127{unit_1_io_out[63]}},unit_1_io_out}; // @[Cordic_HV_Square_Root.scala 185:30]
  wire [190:0] _temp_out_T_3 = $signed(_GEN_0) << u_cnt_1[7:1]; // @[Cordic_HV_Square_Root.scala 185:30]
  wire [190:0] _GEN_2 = $signed(cnt_reg_14) > 8'sh0 ? $signed({{127{_temp_out_T_1[63]}},_temp_out_T_1}) : $signed(
    _temp_out_T_3); // @[Cordic_HV_Square_Root.scala 179:43 182:14 185:14]
  wire [63:0] temp_out = _GEN_2[63:0]; // @[Cordic_HV_Square_Root.scala 155:34]
  wire [63:0] _io_out_T_2 = 64'sh0 - $signed(temp_out); // @[Cordic_HV_Square_Root.scala 191:15]
  shift_range_1_8 unit ( // @[Cordic_HV_Square_Root.scala 130:22]
    .io_x(unit_io_x),
    .io_out(unit_io_out),
    .io_cnt(unit_io_cnt)
  );
  cordic_hv_square_root_origin unit_1 ( // @[Cordic_HV_Square_Root.scala 176:20]
    .clock(unit_1_clock),
    .reset(unit_1_reset),
    .io_in(unit_1_io_in),
    .io_out(unit_1_io_out)
  );
  assign io_out = flag ? $signed(temp_out) : $signed(_io_out_T_2); // @[Cordic_HV_Square_Root.scala 188:14 189:12 191:12]
  assign unit_io_x = flag ? $signed(io_in) : $signed(_temp_in_T_2); // @[Cordic_HV_Square_Root.scala 156:51 157:13 160:13]
  assign unit_1_clock = clock;
  assign unit_1_reset = reset;
  assign unit_1_io_in = unit_io_out; // @[Cordic_HV_Square_Root.scala 177:14]
  always @(posedge clock) begin
    if (reset) begin // @[Cordic_HV_Square_Root.scala 167:35]
      cnt_reg_0 <= 8'sh0; // @[Cordic_HV_Square_Root.scala 167:35]
    end else begin
      cnt_reg_0 <= unit_io_cnt; // @[Cordic_HV_Square_Root.scala 170:18]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 167:35]
      cnt_reg_1 <= 8'sh0; // @[Cordic_HV_Square_Root.scala 167:35]
    end else begin
      cnt_reg_1 <= cnt_reg_0; // @[Cordic_HV_Square_Root.scala 172:18]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 167:35]
      cnt_reg_2 <= 8'sh0; // @[Cordic_HV_Square_Root.scala 167:35]
    end else begin
      cnt_reg_2 <= cnt_reg_1; // @[Cordic_HV_Square_Root.scala 172:18]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 167:35]
      cnt_reg_3 <= 8'sh0; // @[Cordic_HV_Square_Root.scala 167:35]
    end else begin
      cnt_reg_3 <= cnt_reg_2; // @[Cordic_HV_Square_Root.scala 172:18]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 167:35]
      cnt_reg_4 <= 8'sh0; // @[Cordic_HV_Square_Root.scala 167:35]
    end else begin
      cnt_reg_4 <= cnt_reg_3; // @[Cordic_HV_Square_Root.scala 172:18]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 167:35]
      cnt_reg_5 <= 8'sh0; // @[Cordic_HV_Square_Root.scala 167:35]
    end else begin
      cnt_reg_5 <= cnt_reg_4; // @[Cordic_HV_Square_Root.scala 172:18]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 167:35]
      cnt_reg_6 <= 8'sh0; // @[Cordic_HV_Square_Root.scala 167:35]
    end else begin
      cnt_reg_6 <= cnt_reg_5; // @[Cordic_HV_Square_Root.scala 172:18]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 167:35]
      cnt_reg_7 <= 8'sh0; // @[Cordic_HV_Square_Root.scala 167:35]
    end else begin
      cnt_reg_7 <= cnt_reg_6; // @[Cordic_HV_Square_Root.scala 172:18]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 167:35]
      cnt_reg_8 <= 8'sh0; // @[Cordic_HV_Square_Root.scala 167:35]
    end else begin
      cnt_reg_8 <= cnt_reg_7; // @[Cordic_HV_Square_Root.scala 172:18]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 167:35]
      cnt_reg_9 <= 8'sh0; // @[Cordic_HV_Square_Root.scala 167:35]
    end else begin
      cnt_reg_9 <= cnt_reg_8; // @[Cordic_HV_Square_Root.scala 172:18]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 167:35]
      cnt_reg_10 <= 8'sh0; // @[Cordic_HV_Square_Root.scala 167:35]
    end else begin
      cnt_reg_10 <= cnt_reg_9; // @[Cordic_HV_Square_Root.scala 172:18]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 167:35]
      cnt_reg_11 <= 8'sh0; // @[Cordic_HV_Square_Root.scala 167:35]
    end else begin
      cnt_reg_11 <= cnt_reg_10; // @[Cordic_HV_Square_Root.scala 172:18]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 167:35]
      cnt_reg_12 <= 8'sh0; // @[Cordic_HV_Square_Root.scala 167:35]
    end else begin
      cnt_reg_12 <= cnt_reg_11; // @[Cordic_HV_Square_Root.scala 172:18]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 167:35]
      cnt_reg_13 <= 8'sh0; // @[Cordic_HV_Square_Root.scala 167:35]
    end else begin
      cnt_reg_13 <= cnt_reg_12; // @[Cordic_HV_Square_Root.scala 172:18]
    end
    if (reset) begin // @[Cordic_HV_Square_Root.scala 167:35]
      cnt_reg_14 <= 8'sh0; // @[Cordic_HV_Square_Root.scala 167:35]
    end else begin
      cnt_reg_14 <= cnt_reg_13; // @[Cordic_HV_Square_Root.scala 172:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt_reg_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  cnt_reg_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  cnt_reg_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  cnt_reg_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  cnt_reg_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  cnt_reg_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  cnt_reg_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  cnt_reg_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  cnt_reg_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  cnt_reg_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  cnt_reg_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  cnt_reg_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  cnt_reg_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  cnt_reg_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  cnt_reg_14 = _RAND_14[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cordic_complex_square_root(
  input         clock,
  input         reset,
  input  [63:0] io_op_re,
  input  [63:0] io_op_im,
  output [63:0] io_res_re,
  output [63:0] io_res_im
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
`endif // RANDOMIZE_REG_INIT
  wire  io_res_re_unit_clock; // @[Cordic_HV_Square_Root.scala 211:22]
  wire  io_res_re_unit_reset; // @[Cordic_HV_Square_Root.scala 211:22]
  wire [63:0] io_res_re_unit_io_in; // @[Cordic_HV_Square_Root.scala 211:22]
  wire [63:0] io_res_re_unit_io_out; // @[Cordic_HV_Square_Root.scala 211:22]
  wire  io_res_im_unit_clock; // @[Cordic_HV_Square_Root.scala 211:22]
  wire  io_res_im_unit_reset; // @[Cordic_HV_Square_Root.scala 211:22]
  wire [63:0] io_res_im_unit_io_in; // @[Cordic_HV_Square_Root.scala 211:22]
  wire [63:0] io_res_im_unit_io_out; // @[Cordic_HV_Square_Root.scala 211:22]
  reg [63:0] current_x_0; // @[Cordic_Complex_Square_Root.scala 22:43]
  reg [63:0] current_x_1; // @[Cordic_Complex_Square_Root.scala 22:43]
  reg [63:0] current_x_2; // @[Cordic_Complex_Square_Root.scala 22:43]
  reg [63:0] current_x_3; // @[Cordic_Complex_Square_Root.scala 22:43]
  reg [63:0] current_x_4; // @[Cordic_Complex_Square_Root.scala 22:43]
  reg [63:0] current_x_5; // @[Cordic_Complex_Square_Root.scala 22:43]
  reg [63:0] current_x_6; // @[Cordic_Complex_Square_Root.scala 22:43]
  reg [63:0] current_x_7; // @[Cordic_Complex_Square_Root.scala 22:43]
  reg [63:0] current_x_8; // @[Cordic_Complex_Square_Root.scala 22:43]
  reg [63:0] current_x_9; // @[Cordic_Complex_Square_Root.scala 22:43]
  reg [63:0] current_x_10; // @[Cordic_Complex_Square_Root.scala 22:43]
  reg [63:0] current_x_11; // @[Cordic_Complex_Square_Root.scala 22:43]
  reg [63:0] current_x_12; // @[Cordic_Complex_Square_Root.scala 22:43]
  reg [63:0] current_x_13; // @[Cordic_Complex_Square_Root.scala 22:43]
  reg [63:0] current_x_14; // @[Cordic_Complex_Square_Root.scala 22:43]
  reg [63:0] current_y_0; // @[Cordic_Complex_Square_Root.scala 23:43]
  reg [63:0] current_y_1; // @[Cordic_Complex_Square_Root.scala 23:43]
  reg [63:0] current_y_2; // @[Cordic_Complex_Square_Root.scala 23:43]
  reg [63:0] current_y_3; // @[Cordic_Complex_Square_Root.scala 23:43]
  reg [63:0] current_y_4; // @[Cordic_Complex_Square_Root.scala 23:43]
  reg [63:0] current_y_5; // @[Cordic_Complex_Square_Root.scala 23:43]
  reg [63:0] current_y_6; // @[Cordic_Complex_Square_Root.scala 23:43]
  reg [63:0] current_y_7; // @[Cordic_Complex_Square_Root.scala 23:43]
  reg [63:0] current_y_8; // @[Cordic_Complex_Square_Root.scala 23:43]
  reg [63:0] current_y_9; // @[Cordic_Complex_Square_Root.scala 23:43]
  reg [63:0] current_y_10; // @[Cordic_Complex_Square_Root.scala 23:43]
  reg [63:0] current_y_11; // @[Cordic_Complex_Square_Root.scala 23:43]
  reg [63:0] current_y_12; // @[Cordic_Complex_Square_Root.scala 23:43]
  reg [63:0] current_y_13; // @[Cordic_Complex_Square_Root.scala 23:43]
  reg [63:0] reg_x_0; // @[Cordic_Complex_Square_Root.scala 26:39]
  reg [63:0] reg_x_1; // @[Cordic_Complex_Square_Root.scala 26:39]
  reg [63:0] reg_x_2; // @[Cordic_Complex_Square_Root.scala 26:39]
  reg [63:0] reg_x_3; // @[Cordic_Complex_Square_Root.scala 26:39]
  reg [63:0] reg_x_4; // @[Cordic_Complex_Square_Root.scala 26:39]
  reg [63:0] reg_x_5; // @[Cordic_Complex_Square_Root.scala 26:39]
  reg [63:0] reg_x_6; // @[Cordic_Complex_Square_Root.scala 26:39]
  reg [63:0] reg_x_7; // @[Cordic_Complex_Square_Root.scala 26:39]
  reg [63:0] reg_x_8; // @[Cordic_Complex_Square_Root.scala 26:39]
  reg [63:0] reg_x_9; // @[Cordic_Complex_Square_Root.scala 26:39]
  reg [63:0] reg_x_10; // @[Cordic_Complex_Square_Root.scala 26:39]
  reg [63:0] reg_x_11; // @[Cordic_Complex_Square_Root.scala 26:39]
  reg [63:0] reg_x_12; // @[Cordic_Complex_Square_Root.scala 26:39]
  reg [63:0] reg_x_13; // @[Cordic_Complex_Square_Root.scala 26:39]
  reg [63:0] reg_x_14; // @[Cordic_Complex_Square_Root.scala 26:39]
  wire [63:0] _current_x_0_T_3 = $signed(io_op_re) - $signed(io_op_im); // @[Cordic_Complex_Square_Root.scala 36:27]
  wire [63:0] _current_y_0_T_3 = $signed(io_op_im) + $signed(io_op_re); // @[Cordic_Complex_Square_Root.scala 37:27]
  wire [63:0] _current_x_0_T_7 = $signed(io_op_re) + $signed(io_op_im); // @[Cordic_Complex_Square_Root.scala 39:27]
  wire [63:0] _current_y_0_T_7 = $signed(io_op_im) - $signed(io_op_re); // @[Cordic_Complex_Square_Root.scala 40:27]
  wire [62:0] _current_x_1_T = current_y_0[63:1]; // @[Cordic_Complex_Square_Root.scala 45:62]
  wire [63:0] _GEN_30 = {{1{_current_x_1_T[62]}},_current_x_1_T}; // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [63:0] _current_x_1_T_3 = $signed(current_x_0) - $signed(_GEN_30); // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [62:0] _current_y_1_T = current_x_0[63:1]; // @[Cordic_Complex_Square_Root.scala 46:62]
  wire [63:0] _GEN_31 = {{1{_current_y_1_T[62]}},_current_y_1_T}; // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_y_1_T_3 = $signed(current_y_0) + $signed(_GEN_31); // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_x_1_T_7 = $signed(current_x_0) + $signed(_GEN_30); // @[Cordic_Complex_Square_Root.scala 48:42]
  wire [63:0] _current_y_1_T_7 = $signed(current_y_0) - $signed(_GEN_31); // @[Cordic_Complex_Square_Root.scala 49:42]
  wire [61:0] _current_x_2_T = current_y_1[63:2]; // @[Cordic_Complex_Square_Root.scala 45:62]
  wire [63:0] _GEN_34 = {{2{_current_x_2_T[61]}},_current_x_2_T}; // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [63:0] _current_x_2_T_3 = $signed(current_x_1) - $signed(_GEN_34); // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [61:0] _current_y_2_T = current_x_1[63:2]; // @[Cordic_Complex_Square_Root.scala 46:62]
  wire [63:0] _GEN_35 = {{2{_current_y_2_T[61]}},_current_y_2_T}; // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_y_2_T_3 = $signed(current_y_1) + $signed(_GEN_35); // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_x_2_T_7 = $signed(current_x_1) + $signed(_GEN_34); // @[Cordic_Complex_Square_Root.scala 48:42]
  wire [63:0] _current_y_2_T_7 = $signed(current_y_1) - $signed(_GEN_35); // @[Cordic_Complex_Square_Root.scala 49:42]
  wire [60:0] _current_x_3_T = current_y_2[63:3]; // @[Cordic_Complex_Square_Root.scala 45:62]
  wire [63:0] _GEN_38 = {{3{_current_x_3_T[60]}},_current_x_3_T}; // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [63:0] _current_x_3_T_3 = $signed(current_x_2) - $signed(_GEN_38); // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [60:0] _current_y_3_T = current_x_2[63:3]; // @[Cordic_Complex_Square_Root.scala 46:62]
  wire [63:0] _GEN_39 = {{3{_current_y_3_T[60]}},_current_y_3_T}; // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_y_3_T_3 = $signed(current_y_2) + $signed(_GEN_39); // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_x_3_T_7 = $signed(current_x_2) + $signed(_GEN_38); // @[Cordic_Complex_Square_Root.scala 48:42]
  wire [63:0] _current_y_3_T_7 = $signed(current_y_2) - $signed(_GEN_39); // @[Cordic_Complex_Square_Root.scala 49:42]
  wire [59:0] _current_x_4_T = current_y_3[63:4]; // @[Cordic_Complex_Square_Root.scala 45:62]
  wire [63:0] _GEN_42 = {{4{_current_x_4_T[59]}},_current_x_4_T}; // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [63:0] _current_x_4_T_3 = $signed(current_x_3) - $signed(_GEN_42); // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [59:0] _current_y_4_T = current_x_3[63:4]; // @[Cordic_Complex_Square_Root.scala 46:62]
  wire [63:0] _GEN_43 = {{4{_current_y_4_T[59]}},_current_y_4_T}; // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_y_4_T_3 = $signed(current_y_3) + $signed(_GEN_43); // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_x_4_T_7 = $signed(current_x_3) + $signed(_GEN_42); // @[Cordic_Complex_Square_Root.scala 48:42]
  wire [63:0] _current_y_4_T_7 = $signed(current_y_3) - $signed(_GEN_43); // @[Cordic_Complex_Square_Root.scala 49:42]
  wire [58:0] _current_x_5_T = current_y_4[63:5]; // @[Cordic_Complex_Square_Root.scala 45:62]
  wire [63:0] _GEN_46 = {{5{_current_x_5_T[58]}},_current_x_5_T}; // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [63:0] _current_x_5_T_3 = $signed(current_x_4) - $signed(_GEN_46); // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [58:0] _current_y_5_T = current_x_4[63:5]; // @[Cordic_Complex_Square_Root.scala 46:62]
  wire [63:0] _GEN_47 = {{5{_current_y_5_T[58]}},_current_y_5_T}; // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_y_5_T_3 = $signed(current_y_4) + $signed(_GEN_47); // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_x_5_T_7 = $signed(current_x_4) + $signed(_GEN_46); // @[Cordic_Complex_Square_Root.scala 48:42]
  wire [63:0] _current_y_5_T_7 = $signed(current_y_4) - $signed(_GEN_47); // @[Cordic_Complex_Square_Root.scala 49:42]
  wire [57:0] _current_x_6_T = current_y_5[63:6]; // @[Cordic_Complex_Square_Root.scala 45:62]
  wire [63:0] _GEN_50 = {{6{_current_x_6_T[57]}},_current_x_6_T}; // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [63:0] _current_x_6_T_3 = $signed(current_x_5) - $signed(_GEN_50); // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [57:0] _current_y_6_T = current_x_5[63:6]; // @[Cordic_Complex_Square_Root.scala 46:62]
  wire [63:0] _GEN_51 = {{6{_current_y_6_T[57]}},_current_y_6_T}; // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_y_6_T_3 = $signed(current_y_5) + $signed(_GEN_51); // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_x_6_T_7 = $signed(current_x_5) + $signed(_GEN_50); // @[Cordic_Complex_Square_Root.scala 48:42]
  wire [63:0] _current_y_6_T_7 = $signed(current_y_5) - $signed(_GEN_51); // @[Cordic_Complex_Square_Root.scala 49:42]
  wire [56:0] _current_x_7_T = current_y_6[63:7]; // @[Cordic_Complex_Square_Root.scala 45:62]
  wire [63:0] _GEN_54 = {{7{_current_x_7_T[56]}},_current_x_7_T}; // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [63:0] _current_x_7_T_3 = $signed(current_x_6) - $signed(_GEN_54); // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [56:0] _current_y_7_T = current_x_6[63:7]; // @[Cordic_Complex_Square_Root.scala 46:62]
  wire [63:0] _GEN_55 = {{7{_current_y_7_T[56]}},_current_y_7_T}; // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_y_7_T_3 = $signed(current_y_6) + $signed(_GEN_55); // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_x_7_T_7 = $signed(current_x_6) + $signed(_GEN_54); // @[Cordic_Complex_Square_Root.scala 48:42]
  wire [63:0] _current_y_7_T_7 = $signed(current_y_6) - $signed(_GEN_55); // @[Cordic_Complex_Square_Root.scala 49:42]
  wire [55:0] _current_x_8_T = current_y_7[63:8]; // @[Cordic_Complex_Square_Root.scala 45:62]
  wire [63:0] _GEN_58 = {{8{_current_x_8_T[55]}},_current_x_8_T}; // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [63:0] _current_x_8_T_3 = $signed(current_x_7) - $signed(_GEN_58); // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [55:0] _current_y_8_T = current_x_7[63:8]; // @[Cordic_Complex_Square_Root.scala 46:62]
  wire [63:0] _GEN_59 = {{8{_current_y_8_T[55]}},_current_y_8_T}; // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_y_8_T_3 = $signed(current_y_7) + $signed(_GEN_59); // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_x_8_T_7 = $signed(current_x_7) + $signed(_GEN_58); // @[Cordic_Complex_Square_Root.scala 48:42]
  wire [63:0] _current_y_8_T_7 = $signed(current_y_7) - $signed(_GEN_59); // @[Cordic_Complex_Square_Root.scala 49:42]
  wire [54:0] _current_x_9_T = current_y_8[63:9]; // @[Cordic_Complex_Square_Root.scala 45:62]
  wire [63:0] _GEN_62 = {{9{_current_x_9_T[54]}},_current_x_9_T}; // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [63:0] _current_x_9_T_3 = $signed(current_x_8) - $signed(_GEN_62); // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [54:0] _current_y_9_T = current_x_8[63:9]; // @[Cordic_Complex_Square_Root.scala 46:62]
  wire [63:0] _GEN_63 = {{9{_current_y_9_T[54]}},_current_y_9_T}; // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_y_9_T_3 = $signed(current_y_8) + $signed(_GEN_63); // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_x_9_T_7 = $signed(current_x_8) + $signed(_GEN_62); // @[Cordic_Complex_Square_Root.scala 48:42]
  wire [63:0] _current_y_9_T_7 = $signed(current_y_8) - $signed(_GEN_63); // @[Cordic_Complex_Square_Root.scala 49:42]
  wire [53:0] _current_x_10_T = current_y_9[63:10]; // @[Cordic_Complex_Square_Root.scala 45:62]
  wire [63:0] _GEN_66 = {{10{_current_x_10_T[53]}},_current_x_10_T}; // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [63:0] _current_x_10_T_3 = $signed(current_x_9) - $signed(_GEN_66); // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [53:0] _current_y_10_T = current_x_9[63:10]; // @[Cordic_Complex_Square_Root.scala 46:62]
  wire [63:0] _GEN_67 = {{10{_current_y_10_T[53]}},_current_y_10_T}; // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_y_10_T_3 = $signed(current_y_9) + $signed(_GEN_67); // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_x_10_T_7 = $signed(current_x_9) + $signed(_GEN_66); // @[Cordic_Complex_Square_Root.scala 48:42]
  wire [63:0] _current_y_10_T_7 = $signed(current_y_9) - $signed(_GEN_67); // @[Cordic_Complex_Square_Root.scala 49:42]
  wire [52:0] _current_x_11_T = current_y_10[63:11]; // @[Cordic_Complex_Square_Root.scala 45:62]
  wire [63:0] _GEN_70 = {{11{_current_x_11_T[52]}},_current_x_11_T}; // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [63:0] _current_x_11_T_3 = $signed(current_x_10) - $signed(_GEN_70); // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [52:0] _current_y_11_T = current_x_10[63:11]; // @[Cordic_Complex_Square_Root.scala 46:62]
  wire [63:0] _GEN_71 = {{11{_current_y_11_T[52]}},_current_y_11_T}; // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_y_11_T_3 = $signed(current_y_10) + $signed(_GEN_71); // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_x_11_T_7 = $signed(current_x_10) + $signed(_GEN_70); // @[Cordic_Complex_Square_Root.scala 48:42]
  wire [63:0] _current_y_11_T_7 = $signed(current_y_10) - $signed(_GEN_71); // @[Cordic_Complex_Square_Root.scala 49:42]
  wire [51:0] _current_x_12_T = current_y_11[63:12]; // @[Cordic_Complex_Square_Root.scala 45:62]
  wire [63:0] _GEN_74 = {{12{_current_x_12_T[51]}},_current_x_12_T}; // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [63:0] _current_x_12_T_3 = $signed(current_x_11) - $signed(_GEN_74); // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [51:0] _current_y_12_T = current_x_11[63:12]; // @[Cordic_Complex_Square_Root.scala 46:62]
  wire [63:0] _GEN_75 = {{12{_current_y_12_T[51]}},_current_y_12_T}; // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_y_12_T_3 = $signed(current_y_11) + $signed(_GEN_75); // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_x_12_T_7 = $signed(current_x_11) + $signed(_GEN_74); // @[Cordic_Complex_Square_Root.scala 48:42]
  wire [63:0] _current_y_12_T_7 = $signed(current_y_11) - $signed(_GEN_75); // @[Cordic_Complex_Square_Root.scala 49:42]
  wire [50:0] _current_x_13_T = current_y_12[63:13]; // @[Cordic_Complex_Square_Root.scala 45:62]
  wire [63:0] _GEN_78 = {{13{_current_x_13_T[50]}},_current_x_13_T}; // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [63:0] _current_x_13_T_3 = $signed(current_x_12) - $signed(_GEN_78); // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [50:0] _current_y_13_T = current_x_12[63:13]; // @[Cordic_Complex_Square_Root.scala 46:62]
  wire [63:0] _GEN_79 = {{13{_current_y_13_T[50]}},_current_y_13_T}; // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_y_13_T_3 = $signed(current_y_12) + $signed(_GEN_79); // @[Cordic_Complex_Square_Root.scala 46:42]
  wire [63:0] _current_x_13_T_7 = $signed(current_x_12) + $signed(_GEN_78); // @[Cordic_Complex_Square_Root.scala 48:42]
  wire [63:0] _current_y_13_T_7 = $signed(current_y_12) - $signed(_GEN_79); // @[Cordic_Complex_Square_Root.scala 49:42]
  wire [49:0] _current_x_14_T = current_y_13[63:14]; // @[Cordic_Complex_Square_Root.scala 45:62]
  wire [63:0] _GEN_82 = {{14{_current_x_14_T[49]}},_current_x_14_T}; // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [63:0] _current_x_14_T_3 = $signed(current_x_13) - $signed(_GEN_82); // @[Cordic_Complex_Square_Root.scala 45:42]
  wire [63:0] _current_x_14_T_7 = $signed(current_x_13) + $signed(_GEN_82); // @[Cordic_Complex_Square_Root.scala 48:42]
  wire [127:0] temp_cv_out = $signed(current_x_14) * 64'sh9b74eda8; // @[Cordic_Complex_Square_Root.scala 55:50]
  wire [95:0] _GEN_86 = {$signed(reg_x_14), 32'h0}; // @[Cordic_Complex_Square_Root.scala 58:29]
  wire [127:0] _GEN_87 = {{32{_GEN_86[95]}},_GEN_86}; // @[Cordic_Complex_Square_Root.scala 58:29]
  wire [127:0] _next_x_T_2 = $signed(temp_cv_out) + $signed(_GEN_87); // @[Cordic_Complex_Square_Root.scala 58:29]
  wire [126:0] next_x = _next_x_T_2[127:1]; // @[Cordic_Complex_Square_Root.scala 58:58]
  wire [127:0] _next_y_T_2 = $signed(temp_cv_out) - $signed(_GEN_87); // @[Cordic_Complex_Square_Root.scala 59:29]
  wire [126:0] next_y = _next_y_T_2[127:1]; // @[Cordic_Complex_Square_Root.scala 59:58]
  wire [94:0] _GEN_90 = next_x[126:32]; // @[Cordic_HV_Square_Root.scala 212:16]
  wire [94:0] _GEN_92 = next_y[126:32]; // @[Cordic_HV_Square_Root.scala 212:16]
  cordic_hv_square_root io_res_re_unit ( // @[Cordic_HV_Square_Root.scala 211:22]
    .clock(io_res_re_unit_clock),
    .reset(io_res_re_unit_reset),
    .io_in(io_res_re_unit_io_in),
    .io_out(io_res_re_unit_io_out)
  );
  cordic_hv_square_root io_res_im_unit ( // @[Cordic_HV_Square_Root.scala 211:22]
    .clock(io_res_im_unit_clock),
    .reset(io_res_im_unit_reset),
    .io_in(io_res_im_unit_io_in),
    .io_out(io_res_im_unit_io_out)
  );
  assign io_res_re = io_res_re_unit_io_out; // @[Cordic_Complex_Square_Root.scala 60:13]
  assign io_res_im = io_res_im_unit_io_out; // @[Cordic_Complex_Square_Root.scala 61:13]
  assign io_res_re_unit_clock = clock;
  assign io_res_re_unit_reset = reset;
  assign io_res_re_unit_io_in = _GEN_90[63:0]; // @[Cordic_HV_Square_Root.scala 212:16]
  assign io_res_im_unit_clock = clock;
  assign io_res_im_unit_reset = reset;
  assign io_res_im_unit_io_in = _GEN_92[63:0]; // @[Cordic_HV_Square_Root.scala 212:16]
  always @(posedge clock) begin
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 22:43]
      current_x_0 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 22:43]
    end else if ($signed(io_op_im) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 35:73]
      current_x_0 <= _current_x_0_T_3; // @[Cordic_Complex_Square_Root.scala 36:22]
    end else begin
      current_x_0 <= _current_x_0_T_7; // @[Cordic_Complex_Square_Root.scala 39:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 22:43]
      current_x_1 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 22:43]
    end else if ($signed(current_y_0) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_x_1 <= _current_x_1_T_3; // @[Cordic_Complex_Square_Root.scala 45:22]
    end else begin
      current_x_1 <= _current_x_1_T_7; // @[Cordic_Complex_Square_Root.scala 48:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 22:43]
      current_x_2 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 22:43]
    end else if ($signed(current_y_1) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_x_2 <= _current_x_2_T_3; // @[Cordic_Complex_Square_Root.scala 45:22]
    end else begin
      current_x_2 <= _current_x_2_T_7; // @[Cordic_Complex_Square_Root.scala 48:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 22:43]
      current_x_3 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 22:43]
    end else if ($signed(current_y_2) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_x_3 <= _current_x_3_T_3; // @[Cordic_Complex_Square_Root.scala 45:22]
    end else begin
      current_x_3 <= _current_x_3_T_7; // @[Cordic_Complex_Square_Root.scala 48:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 22:43]
      current_x_4 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 22:43]
    end else if ($signed(current_y_3) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_x_4 <= _current_x_4_T_3; // @[Cordic_Complex_Square_Root.scala 45:22]
    end else begin
      current_x_4 <= _current_x_4_T_7; // @[Cordic_Complex_Square_Root.scala 48:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 22:43]
      current_x_5 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 22:43]
    end else if ($signed(current_y_4) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_x_5 <= _current_x_5_T_3; // @[Cordic_Complex_Square_Root.scala 45:22]
    end else begin
      current_x_5 <= _current_x_5_T_7; // @[Cordic_Complex_Square_Root.scala 48:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 22:43]
      current_x_6 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 22:43]
    end else if ($signed(current_y_5) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_x_6 <= _current_x_6_T_3; // @[Cordic_Complex_Square_Root.scala 45:22]
    end else begin
      current_x_6 <= _current_x_6_T_7; // @[Cordic_Complex_Square_Root.scala 48:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 22:43]
      current_x_7 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 22:43]
    end else if ($signed(current_y_6) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_x_7 <= _current_x_7_T_3; // @[Cordic_Complex_Square_Root.scala 45:22]
    end else begin
      current_x_7 <= _current_x_7_T_7; // @[Cordic_Complex_Square_Root.scala 48:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 22:43]
      current_x_8 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 22:43]
    end else if ($signed(current_y_7) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_x_8 <= _current_x_8_T_3; // @[Cordic_Complex_Square_Root.scala 45:22]
    end else begin
      current_x_8 <= _current_x_8_T_7; // @[Cordic_Complex_Square_Root.scala 48:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 22:43]
      current_x_9 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 22:43]
    end else if ($signed(current_y_8) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_x_9 <= _current_x_9_T_3; // @[Cordic_Complex_Square_Root.scala 45:22]
    end else begin
      current_x_9 <= _current_x_9_T_7; // @[Cordic_Complex_Square_Root.scala 48:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 22:43]
      current_x_10 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 22:43]
    end else if ($signed(current_y_9) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_x_10 <= _current_x_10_T_3; // @[Cordic_Complex_Square_Root.scala 45:22]
    end else begin
      current_x_10 <= _current_x_10_T_7; // @[Cordic_Complex_Square_Root.scala 48:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 22:43]
      current_x_11 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 22:43]
    end else if ($signed(current_y_10) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_x_11 <= _current_x_11_T_3; // @[Cordic_Complex_Square_Root.scala 45:22]
    end else begin
      current_x_11 <= _current_x_11_T_7; // @[Cordic_Complex_Square_Root.scala 48:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 22:43]
      current_x_12 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 22:43]
    end else if ($signed(current_y_11) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_x_12 <= _current_x_12_T_3; // @[Cordic_Complex_Square_Root.scala 45:22]
    end else begin
      current_x_12 <= _current_x_12_T_7; // @[Cordic_Complex_Square_Root.scala 48:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 22:43]
      current_x_13 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 22:43]
    end else if ($signed(current_y_12) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_x_13 <= _current_x_13_T_3; // @[Cordic_Complex_Square_Root.scala 45:22]
    end else begin
      current_x_13 <= _current_x_13_T_7; // @[Cordic_Complex_Square_Root.scala 48:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 22:43]
      current_x_14 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 22:43]
    end else if ($signed(current_y_13) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_x_14 <= _current_x_14_T_3; // @[Cordic_Complex_Square_Root.scala 45:22]
    end else begin
      current_x_14 <= _current_x_14_T_7; // @[Cordic_Complex_Square_Root.scala 48:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 23:43]
      current_y_0 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 23:43]
    end else if ($signed(io_op_im) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 35:73]
      current_y_0 <= _current_y_0_T_3; // @[Cordic_Complex_Square_Root.scala 37:22]
    end else begin
      current_y_0 <= _current_y_0_T_7; // @[Cordic_Complex_Square_Root.scala 40:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 23:43]
      current_y_1 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 23:43]
    end else if ($signed(current_y_0) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_y_1 <= _current_y_1_T_3; // @[Cordic_Complex_Square_Root.scala 46:22]
    end else begin
      current_y_1 <= _current_y_1_T_7; // @[Cordic_Complex_Square_Root.scala 49:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 23:43]
      current_y_2 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 23:43]
    end else if ($signed(current_y_1) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_y_2 <= _current_y_2_T_3; // @[Cordic_Complex_Square_Root.scala 46:22]
    end else begin
      current_y_2 <= _current_y_2_T_7; // @[Cordic_Complex_Square_Root.scala 49:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 23:43]
      current_y_3 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 23:43]
    end else if ($signed(current_y_2) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_y_3 <= _current_y_3_T_3; // @[Cordic_Complex_Square_Root.scala 46:22]
    end else begin
      current_y_3 <= _current_y_3_T_7; // @[Cordic_Complex_Square_Root.scala 49:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 23:43]
      current_y_4 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 23:43]
    end else if ($signed(current_y_3) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_y_4 <= _current_y_4_T_3; // @[Cordic_Complex_Square_Root.scala 46:22]
    end else begin
      current_y_4 <= _current_y_4_T_7; // @[Cordic_Complex_Square_Root.scala 49:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 23:43]
      current_y_5 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 23:43]
    end else if ($signed(current_y_4) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_y_5 <= _current_y_5_T_3; // @[Cordic_Complex_Square_Root.scala 46:22]
    end else begin
      current_y_5 <= _current_y_5_T_7; // @[Cordic_Complex_Square_Root.scala 49:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 23:43]
      current_y_6 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 23:43]
    end else if ($signed(current_y_5) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_y_6 <= _current_y_6_T_3; // @[Cordic_Complex_Square_Root.scala 46:22]
    end else begin
      current_y_6 <= _current_y_6_T_7; // @[Cordic_Complex_Square_Root.scala 49:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 23:43]
      current_y_7 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 23:43]
    end else if ($signed(current_y_6) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_y_7 <= _current_y_7_T_3; // @[Cordic_Complex_Square_Root.scala 46:22]
    end else begin
      current_y_7 <= _current_y_7_T_7; // @[Cordic_Complex_Square_Root.scala 49:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 23:43]
      current_y_8 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 23:43]
    end else if ($signed(current_y_7) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_y_8 <= _current_y_8_T_3; // @[Cordic_Complex_Square_Root.scala 46:22]
    end else begin
      current_y_8 <= _current_y_8_T_7; // @[Cordic_Complex_Square_Root.scala 49:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 23:43]
      current_y_9 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 23:43]
    end else if ($signed(current_y_8) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_y_9 <= _current_y_9_T_3; // @[Cordic_Complex_Square_Root.scala 46:22]
    end else begin
      current_y_9 <= _current_y_9_T_7; // @[Cordic_Complex_Square_Root.scala 49:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 23:43]
      current_y_10 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 23:43]
    end else if ($signed(current_y_9) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_y_10 <= _current_y_10_T_3; // @[Cordic_Complex_Square_Root.scala 46:22]
    end else begin
      current_y_10 <= _current_y_10_T_7; // @[Cordic_Complex_Square_Root.scala 49:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 23:43]
      current_y_11 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 23:43]
    end else if ($signed(current_y_10) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_y_11 <= _current_y_11_T_3; // @[Cordic_Complex_Square_Root.scala 46:22]
    end else begin
      current_y_11 <= _current_y_11_T_7; // @[Cordic_Complex_Square_Root.scala 49:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 23:43]
      current_y_12 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 23:43]
    end else if ($signed(current_y_11) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_y_12 <= _current_y_12_T_3; // @[Cordic_Complex_Square_Root.scala 46:22]
    end else begin
      current_y_12 <= _current_y_12_T_7; // @[Cordic_Complex_Square_Root.scala 49:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 23:43]
      current_y_13 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 23:43]
    end else if ($signed(current_y_12) < 64'sh0) begin // @[Cordic_Complex_Square_Root.scala 44:88]
      current_y_13 <= _current_y_13_T_3; // @[Cordic_Complex_Square_Root.scala 46:22]
    end else begin
      current_y_13 <= _current_y_13_T_7; // @[Cordic_Complex_Square_Root.scala 49:22]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 26:39]
      reg_x_0 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 26:39]
    end else begin
      reg_x_0 <= io_op_re; // @[Cordic_Complex_Square_Root.scala 33:16]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 26:39]
      reg_x_1 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 26:39]
    end else begin
      reg_x_1 <= reg_x_0; // @[Cordic_Complex_Square_Root.scala 43:16]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 26:39]
      reg_x_2 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 26:39]
    end else begin
      reg_x_2 <= reg_x_1; // @[Cordic_Complex_Square_Root.scala 43:16]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 26:39]
      reg_x_3 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 26:39]
    end else begin
      reg_x_3 <= reg_x_2; // @[Cordic_Complex_Square_Root.scala 43:16]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 26:39]
      reg_x_4 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 26:39]
    end else begin
      reg_x_4 <= reg_x_3; // @[Cordic_Complex_Square_Root.scala 43:16]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 26:39]
      reg_x_5 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 26:39]
    end else begin
      reg_x_5 <= reg_x_4; // @[Cordic_Complex_Square_Root.scala 43:16]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 26:39]
      reg_x_6 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 26:39]
    end else begin
      reg_x_6 <= reg_x_5; // @[Cordic_Complex_Square_Root.scala 43:16]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 26:39]
      reg_x_7 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 26:39]
    end else begin
      reg_x_7 <= reg_x_6; // @[Cordic_Complex_Square_Root.scala 43:16]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 26:39]
      reg_x_8 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 26:39]
    end else begin
      reg_x_8 <= reg_x_7; // @[Cordic_Complex_Square_Root.scala 43:16]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 26:39]
      reg_x_9 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 26:39]
    end else begin
      reg_x_9 <= reg_x_8; // @[Cordic_Complex_Square_Root.scala 43:16]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 26:39]
      reg_x_10 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 26:39]
    end else begin
      reg_x_10 <= reg_x_9; // @[Cordic_Complex_Square_Root.scala 43:16]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 26:39]
      reg_x_11 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 26:39]
    end else begin
      reg_x_11 <= reg_x_10; // @[Cordic_Complex_Square_Root.scala 43:16]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 26:39]
      reg_x_12 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 26:39]
    end else begin
      reg_x_12 <= reg_x_11; // @[Cordic_Complex_Square_Root.scala 43:16]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 26:39]
      reg_x_13 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 26:39]
    end else begin
      reg_x_13 <= reg_x_12; // @[Cordic_Complex_Square_Root.scala 43:16]
    end
    if (reset) begin // @[Cordic_Complex_Square_Root.scala 26:39]
      reg_x_14 <= 64'sh0; // @[Cordic_Complex_Square_Root.scala 26:39]
    end else begin
      reg_x_14 <= reg_x_13; // @[Cordic_Complex_Square_Root.scala 43:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  current_x_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  current_x_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  current_x_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  current_x_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  current_x_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  current_x_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  current_x_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  current_x_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  current_x_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  current_x_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  current_x_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  current_x_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  current_x_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  current_x_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  current_x_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  current_y_0 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  current_y_1 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  current_y_2 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  current_y_3 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  current_y_4 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  current_y_5 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  current_y_6 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  current_y_7 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  current_y_8 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  current_y_9 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  current_y_10 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  current_y_11 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  current_y_12 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  current_y_13 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  reg_x_0 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  reg_x_1 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  reg_x_2 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  reg_x_3 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  reg_x_4 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  reg_x_5 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  reg_x_6 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  reg_x_7 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  reg_x_8 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  reg_x_9 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  reg_x_10 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  reg_x_11 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  reg_x_12 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  reg_x_13 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  reg_x_14 = _RAND_43[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CORDIC_CV_ORIGIN(
  input         clock,
  input         reset,
  input  [63:0] io_x,
  input  [63:0] io_y,
  output [63:0] io_theta,
  output [63:0] io_r
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] current_x_0; // @[Cordic_CV.scala 40:43]
  reg [63:0] current_x_1; // @[Cordic_CV.scala 40:43]
  reg [63:0] current_x_2; // @[Cordic_CV.scala 40:43]
  reg [63:0] current_x_3; // @[Cordic_CV.scala 40:43]
  reg [63:0] current_x_4; // @[Cordic_CV.scala 40:43]
  reg [63:0] current_x_5; // @[Cordic_CV.scala 40:43]
  reg [63:0] current_x_6; // @[Cordic_CV.scala 40:43]
  reg [63:0] current_x_7; // @[Cordic_CV.scala 40:43]
  reg [63:0] current_x_8; // @[Cordic_CV.scala 40:43]
  reg [63:0] current_x_9; // @[Cordic_CV.scala 40:43]
  reg [63:0] current_x_10; // @[Cordic_CV.scala 40:43]
  reg [63:0] current_x_11; // @[Cordic_CV.scala 40:43]
  reg [63:0] current_x_12; // @[Cordic_CV.scala 40:43]
  reg [63:0] current_x_13; // @[Cordic_CV.scala 40:43]
  reg [63:0] current_x_14; // @[Cordic_CV.scala 40:43]
  reg [63:0] current_y_0; // @[Cordic_CV.scala 41:43]
  reg [63:0] current_y_1; // @[Cordic_CV.scala 41:43]
  reg [63:0] current_y_2; // @[Cordic_CV.scala 41:43]
  reg [63:0] current_y_3; // @[Cordic_CV.scala 41:43]
  reg [63:0] current_y_4; // @[Cordic_CV.scala 41:43]
  reg [63:0] current_y_5; // @[Cordic_CV.scala 41:43]
  reg [63:0] current_y_6; // @[Cordic_CV.scala 41:43]
  reg [63:0] current_y_7; // @[Cordic_CV.scala 41:43]
  reg [63:0] current_y_8; // @[Cordic_CV.scala 41:43]
  reg [63:0] current_y_9; // @[Cordic_CV.scala 41:43]
  reg [63:0] current_y_10; // @[Cordic_CV.scala 41:43]
  reg [63:0] current_y_11; // @[Cordic_CV.scala 41:43]
  reg [63:0] current_y_12; // @[Cordic_CV.scala 41:43]
  reg [63:0] current_y_13; // @[Cordic_CV.scala 41:43]
  reg [63:0] current_theta_0; // @[Cordic_CV.scala 42:47]
  reg [63:0] current_theta_1; // @[Cordic_CV.scala 42:47]
  reg [63:0] current_theta_2; // @[Cordic_CV.scala 42:47]
  reg [63:0] current_theta_3; // @[Cordic_CV.scala 42:47]
  reg [63:0] current_theta_4; // @[Cordic_CV.scala 42:47]
  reg [63:0] current_theta_5; // @[Cordic_CV.scala 42:47]
  reg [63:0] current_theta_6; // @[Cordic_CV.scala 42:47]
  reg [63:0] current_theta_7; // @[Cordic_CV.scala 42:47]
  reg [63:0] current_theta_8; // @[Cordic_CV.scala 42:47]
  reg [63:0] current_theta_9; // @[Cordic_CV.scala 42:47]
  reg [63:0] current_theta_10; // @[Cordic_CV.scala 42:47]
  reg [63:0] current_theta_11; // @[Cordic_CV.scala 42:47]
  reg [63:0] current_theta_12; // @[Cordic_CV.scala 42:47]
  reg [63:0] current_theta_13; // @[Cordic_CV.scala 42:47]
  reg [63:0] current_theta_14; // @[Cordic_CV.scala 42:47]
  wire [63:0] _current_x_0_T_3 = $signed(io_x) - $signed(io_y); // @[Cordic_CV.scala 52:30]
  wire [63:0] _current_y_0_T_3 = $signed(io_y) + $signed(io_x); // @[Cordic_CV.scala 53:30]
  wire [63:0] _current_theta_0_T_2 = 64'sh0 - 64'sh2d00000000; // @[Cordic_CV.scala 54:29]
  wire [63:0] _current_x_0_T_7 = $signed(io_x) + $signed(io_y); // @[Cordic_CV.scala 56:30]
  wire [63:0] _current_y_0_T_7 = $signed(io_y) - $signed(io_x); // @[Cordic_CV.scala 57:30]
  wire [62:0] _current_x_1_T = current_y_0[63:1]; // @[Cordic_CV.scala 62:62]
  wire [63:0] _GEN_45 = {{1{_current_x_1_T[62]}},_current_x_1_T}; // @[Cordic_CV.scala 62:42]
  wire [63:0] _current_x_1_T_3 = $signed(current_x_0) - $signed(_GEN_45); // @[Cordic_CV.scala 62:42]
  wire [62:0] _current_y_1_T = current_x_0[63:1]; // @[Cordic_CV.scala 63:62]
  wire [63:0] _GEN_46 = {{1{_current_y_1_T[62]}},_current_y_1_T}; // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_y_1_T_3 = $signed(current_y_0) + $signed(_GEN_46); // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_theta_1_T_2 = $signed(current_theta_0) - 64'sh1a90a731a6; // @[Cordic_CV.scala 64:50]
  wire [63:0] _current_x_1_T_7 = $signed(current_x_0) + $signed(_GEN_45); // @[Cordic_CV.scala 66:42]
  wire [63:0] _current_y_1_T_7 = $signed(current_y_0) - $signed(_GEN_46); // @[Cordic_CV.scala 67:42]
  wire [63:0] _current_theta_1_T_5 = $signed(current_theta_0) + 64'sh1a90a731a6; // @[Cordic_CV.scala 68:50]
  wire [61:0] _current_x_2_T = current_y_1[63:2]; // @[Cordic_CV.scala 62:62]
  wire [63:0] _GEN_49 = {{2{_current_x_2_T[61]}},_current_x_2_T}; // @[Cordic_CV.scala 62:42]
  wire [63:0] _current_x_2_T_3 = $signed(current_x_1) - $signed(_GEN_49); // @[Cordic_CV.scala 62:42]
  wire [61:0] _current_y_2_T = current_x_1[63:2]; // @[Cordic_CV.scala 63:62]
  wire [63:0] _GEN_50 = {{2{_current_y_2_T[61]}},_current_y_2_T}; // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_y_2_T_3 = $signed(current_y_1) + $signed(_GEN_50); // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_theta_2_T_2 = $signed(current_theta_1) - 64'she0947407d; // @[Cordic_CV.scala 64:50]
  wire [63:0] _current_x_2_T_7 = $signed(current_x_1) + $signed(_GEN_49); // @[Cordic_CV.scala 66:42]
  wire [63:0] _current_y_2_T_7 = $signed(current_y_1) - $signed(_GEN_50); // @[Cordic_CV.scala 67:42]
  wire [63:0] _current_theta_2_T_5 = $signed(current_theta_1) + 64'she0947407d; // @[Cordic_CV.scala 68:50]
  wire [60:0] _current_x_3_T = current_y_2[63:3]; // @[Cordic_CV.scala 62:62]
  wire [63:0] _GEN_53 = {{3{_current_x_3_T[60]}},_current_x_3_T}; // @[Cordic_CV.scala 62:42]
  wire [63:0] _current_x_3_T_3 = $signed(current_x_2) - $signed(_GEN_53); // @[Cordic_CV.scala 62:42]
  wire [60:0] _current_y_3_T = current_x_2[63:3]; // @[Cordic_CV.scala 63:62]
  wire [63:0] _GEN_54 = {{3{_current_y_3_T[60]}},_current_y_3_T}; // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_y_3_T_3 = $signed(current_y_2) + $signed(_GEN_54); // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_theta_3_T_2 = $signed(current_theta_2) - 64'sh72001124a; // @[Cordic_CV.scala 64:50]
  wire [63:0] _current_x_3_T_7 = $signed(current_x_2) + $signed(_GEN_53); // @[Cordic_CV.scala 66:42]
  wire [63:0] _current_y_3_T_7 = $signed(current_y_2) - $signed(_GEN_54); // @[Cordic_CV.scala 67:42]
  wire [63:0] _current_theta_3_T_5 = $signed(current_theta_2) + 64'sh72001124a; // @[Cordic_CV.scala 68:50]
  wire [59:0] _current_x_4_T = current_y_3[63:4]; // @[Cordic_CV.scala 62:62]
  wire [63:0] _GEN_57 = {{4{_current_x_4_T[59]}},_current_x_4_T}; // @[Cordic_CV.scala 62:42]
  wire [63:0] _current_x_4_T_3 = $signed(current_x_3) - $signed(_GEN_57); // @[Cordic_CV.scala 62:42]
  wire [59:0] _current_y_4_T = current_x_3[63:4]; // @[Cordic_CV.scala 63:62]
  wire [63:0] _GEN_58 = {{4{_current_y_4_T[59]}},_current_y_4_T}; // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_y_4_T_3 = $signed(current_y_3) + $signed(_GEN_58); // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_theta_4_T_2 = $signed(current_theta_3) - 64'sh3938aa64c; // @[Cordic_CV.scala 64:50]
  wire [63:0] _current_x_4_T_7 = $signed(current_x_3) + $signed(_GEN_57); // @[Cordic_CV.scala 66:42]
  wire [63:0] _current_y_4_T_7 = $signed(current_y_3) - $signed(_GEN_58); // @[Cordic_CV.scala 67:42]
  wire [63:0] _current_theta_4_T_5 = $signed(current_theta_3) + 64'sh3938aa64c; // @[Cordic_CV.scala 68:50]
  wire [58:0] _current_x_5_T = current_y_4[63:5]; // @[Cordic_CV.scala 62:62]
  wire [63:0] _GEN_61 = {{5{_current_x_5_T[58]}},_current_x_5_T}; // @[Cordic_CV.scala 62:42]
  wire [63:0] _current_x_5_T_3 = $signed(current_x_4) - $signed(_GEN_61); // @[Cordic_CV.scala 62:42]
  wire [58:0] _current_y_5_T = current_x_4[63:5]; // @[Cordic_CV.scala 63:62]
  wire [63:0] _GEN_62 = {{5{_current_y_5_T[58]}},_current_y_5_T}; // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_y_5_T_3 = $signed(current_y_4) + $signed(_GEN_62); // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_theta_5_T_2 = $signed(current_theta_4) - 64'sh1ca3794e5; // @[Cordic_CV.scala 64:50]
  wire [63:0] _current_x_5_T_7 = $signed(current_x_4) + $signed(_GEN_61); // @[Cordic_CV.scala 66:42]
  wire [63:0] _current_y_5_T_7 = $signed(current_y_4) - $signed(_GEN_62); // @[Cordic_CV.scala 67:42]
  wire [63:0] _current_theta_5_T_5 = $signed(current_theta_4) + 64'sh1ca3794e5; // @[Cordic_CV.scala 68:50]
  wire [57:0] _current_x_6_T = current_y_5[63:6]; // @[Cordic_CV.scala 62:62]
  wire [63:0] _GEN_65 = {{6{_current_x_6_T[57]}},_current_x_6_T}; // @[Cordic_CV.scala 62:42]
  wire [63:0] _current_x_6_T_3 = $signed(current_x_5) - $signed(_GEN_65); // @[Cordic_CV.scala 62:42]
  wire [57:0] _current_y_6_T = current_x_5[63:6]; // @[Cordic_CV.scala 63:62]
  wire [63:0] _GEN_66 = {{6{_current_y_6_T[57]}},_current_y_6_T}; // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_y_6_T_3 = $signed(current_y_5) + $signed(_GEN_66); // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_theta_6_T_2 = $signed(current_theta_5) - 64'she52a1ab2; // @[Cordic_CV.scala 64:50]
  wire [63:0] _current_x_6_T_7 = $signed(current_x_5) + $signed(_GEN_65); // @[Cordic_CV.scala 66:42]
  wire [63:0] _current_y_6_T_7 = $signed(current_y_5) - $signed(_GEN_66); // @[Cordic_CV.scala 67:42]
  wire [63:0] _current_theta_6_T_5 = $signed(current_theta_5) + 64'she52a1ab2; // @[Cordic_CV.scala 68:50]
  wire [56:0] _current_x_7_T = current_y_6[63:7]; // @[Cordic_CV.scala 62:62]
  wire [63:0] _GEN_69 = {{7{_current_x_7_T[56]}},_current_x_7_T}; // @[Cordic_CV.scala 62:42]
  wire [63:0] _current_x_7_T_3 = $signed(current_x_6) - $signed(_GEN_69); // @[Cordic_CV.scala 62:42]
  wire [56:0] _current_y_7_T = current_x_6[63:7]; // @[Cordic_CV.scala 63:62]
  wire [63:0] _GEN_70 = {{7{_current_y_7_T[56]}},_current_y_7_T}; // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_y_7_T_3 = $signed(current_y_6) + $signed(_GEN_70); // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_theta_7_T_2 = $signed(current_theta_6) - 64'sh7296d7a1; // @[Cordic_CV.scala 64:50]
  wire [63:0] _current_x_7_T_7 = $signed(current_x_6) + $signed(_GEN_69); // @[Cordic_CV.scala 66:42]
  wire [63:0] _current_y_7_T_7 = $signed(current_y_6) - $signed(_GEN_70); // @[Cordic_CV.scala 67:42]
  wire [63:0] _current_theta_7_T_5 = $signed(current_theta_6) + 64'sh7296d7a1; // @[Cordic_CV.scala 68:50]
  wire [55:0] _current_x_8_T = current_y_7[63:8]; // @[Cordic_CV.scala 62:62]
  wire [63:0] _GEN_73 = {{8{_current_x_8_T[55]}},_current_x_8_T}; // @[Cordic_CV.scala 62:42]
  wire [63:0] _current_x_8_T_3 = $signed(current_x_7) - $signed(_GEN_73); // @[Cordic_CV.scala 62:42]
  wire [55:0] _current_y_8_T = current_x_7[63:8]; // @[Cordic_CV.scala 63:62]
  wire [63:0] _GEN_74 = {{8{_current_y_8_T[55]}},_current_y_8_T}; // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_y_8_T_3 = $signed(current_y_7) + $signed(_GEN_74); // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_theta_8_T_2 = $signed(current_theta_7) - 64'sh394ba51c; // @[Cordic_CV.scala 64:50]
  wire [63:0] _current_x_8_T_7 = $signed(current_x_7) + $signed(_GEN_73); // @[Cordic_CV.scala 66:42]
  wire [63:0] _current_y_8_T_7 = $signed(current_y_7) - $signed(_GEN_74); // @[Cordic_CV.scala 67:42]
  wire [63:0] _current_theta_8_T_5 = $signed(current_theta_7) + 64'sh394ba51c; // @[Cordic_CV.scala 68:50]
  wire [54:0] _current_x_9_T = current_y_8[63:9]; // @[Cordic_CV.scala 62:62]
  wire [63:0] _GEN_77 = {{9{_current_x_9_T[54]}},_current_x_9_T}; // @[Cordic_CV.scala 62:42]
  wire [63:0] _current_x_9_T_3 = $signed(current_x_8) - $signed(_GEN_77); // @[Cordic_CV.scala 62:42]
  wire [54:0] _current_y_9_T = current_x_8[63:9]; // @[Cordic_CV.scala 63:62]
  wire [63:0] _GEN_78 = {{9{_current_y_9_T[54]}},_current_y_9_T}; // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_y_9_T_3 = $signed(current_y_8) + $signed(_GEN_78); // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_theta_9_T_2 = $signed(current_theta_8) - 64'sh1ca5d9b7; // @[Cordic_CV.scala 64:50]
  wire [63:0] _current_x_9_T_7 = $signed(current_x_8) + $signed(_GEN_77); // @[Cordic_CV.scala 66:42]
  wire [63:0] _current_y_9_T_7 = $signed(current_y_8) - $signed(_GEN_78); // @[Cordic_CV.scala 67:42]
  wire [63:0] _current_theta_9_T_5 = $signed(current_theta_8) + 64'sh1ca5d9b7; // @[Cordic_CV.scala 68:50]
  wire [53:0] _current_x_10_T = current_y_9[63:10]; // @[Cordic_CV.scala 62:62]
  wire [63:0] _GEN_81 = {{10{_current_x_10_T[53]}},_current_x_10_T}; // @[Cordic_CV.scala 62:42]
  wire [63:0] _current_x_10_T_3 = $signed(current_x_9) - $signed(_GEN_81); // @[Cordic_CV.scala 62:42]
  wire [53:0] _current_y_10_T = current_x_9[63:10]; // @[Cordic_CV.scala 63:62]
  wire [63:0] _GEN_82 = {{10{_current_y_10_T[53]}},_current_y_10_T}; // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_y_10_T_3 = $signed(current_y_9) + $signed(_GEN_82); // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_theta_10_T_2 = $signed(current_theta_9) - 64'she52edc1; // @[Cordic_CV.scala 64:50]
  wire [63:0] _current_x_10_T_7 = $signed(current_x_9) + $signed(_GEN_81); // @[Cordic_CV.scala 66:42]
  wire [63:0] _current_y_10_T_7 = $signed(current_y_9) - $signed(_GEN_82); // @[Cordic_CV.scala 67:42]
  wire [63:0] _current_theta_10_T_5 = $signed(current_theta_9) + 64'she52edc1; // @[Cordic_CV.scala 68:50]
  wire [52:0] _current_x_11_T = current_y_10[63:11]; // @[Cordic_CV.scala 62:62]
  wire [63:0] _GEN_85 = {{11{_current_x_11_T[52]}},_current_x_11_T}; // @[Cordic_CV.scala 62:42]
  wire [63:0] _current_x_11_T_3 = $signed(current_x_10) - $signed(_GEN_85); // @[Cordic_CV.scala 62:42]
  wire [52:0] _current_y_11_T = current_x_10[63:11]; // @[Cordic_CV.scala 63:62]
  wire [63:0] _GEN_86 = {{11{_current_y_11_T[52]}},_current_y_11_T}; // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_y_11_T_3 = $signed(current_y_10) + $signed(_GEN_86); // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_theta_11_T_2 = $signed(current_theta_10) - 64'sh72976fd; // @[Cordic_CV.scala 64:50]
  wire [63:0] _current_x_11_T_7 = $signed(current_x_10) + $signed(_GEN_85); // @[Cordic_CV.scala 66:42]
  wire [63:0] _current_y_11_T_7 = $signed(current_y_10) - $signed(_GEN_86); // @[Cordic_CV.scala 67:42]
  wire [63:0] _current_theta_11_T_5 = $signed(current_theta_10) + 64'sh72976fd; // @[Cordic_CV.scala 68:50]
  wire [51:0] _current_x_12_T = current_y_11[63:12]; // @[Cordic_CV.scala 62:62]
  wire [63:0] _GEN_89 = {{12{_current_x_12_T[51]}},_current_x_12_T}; // @[Cordic_CV.scala 62:42]
  wire [63:0] _current_x_12_T_3 = $signed(current_x_11) - $signed(_GEN_89); // @[Cordic_CV.scala 62:42]
  wire [51:0] _current_y_12_T = current_x_11[63:12]; // @[Cordic_CV.scala 63:62]
  wire [63:0] _GEN_90 = {{12{_current_y_12_T[51]}},_current_y_12_T}; // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_y_12_T_3 = $signed(current_y_11) + $signed(_GEN_90); // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_theta_12_T_2 = $signed(current_theta_11) - 64'sh394bb82; // @[Cordic_CV.scala 64:50]
  wire [63:0] _current_x_12_T_7 = $signed(current_x_11) + $signed(_GEN_89); // @[Cordic_CV.scala 66:42]
  wire [63:0] _current_y_12_T_7 = $signed(current_y_11) - $signed(_GEN_90); // @[Cordic_CV.scala 67:42]
  wire [63:0] _current_theta_12_T_5 = $signed(current_theta_11) + 64'sh394bb82; // @[Cordic_CV.scala 68:50]
  wire [50:0] _current_x_13_T = current_y_12[63:13]; // @[Cordic_CV.scala 62:62]
  wire [63:0] _GEN_93 = {{13{_current_x_13_T[50]}},_current_x_13_T}; // @[Cordic_CV.scala 62:42]
  wire [63:0] _current_x_13_T_3 = $signed(current_x_12) - $signed(_GEN_93); // @[Cordic_CV.scala 62:42]
  wire [50:0] _current_y_13_T = current_x_12[63:13]; // @[Cordic_CV.scala 63:62]
  wire [63:0] _GEN_94 = {{13{_current_y_13_T[50]}},_current_y_13_T}; // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_y_13_T_3 = $signed(current_y_12) + $signed(_GEN_94); // @[Cordic_CV.scala 63:42]
  wire [63:0] _current_theta_13_T_2 = $signed(current_theta_12) - 64'sh1ca5dc2; // @[Cordic_CV.scala 64:50]
  wire [63:0] _current_x_13_T_7 = $signed(current_x_12) + $signed(_GEN_93); // @[Cordic_CV.scala 66:42]
  wire [63:0] _current_y_13_T_7 = $signed(current_y_12) - $signed(_GEN_94); // @[Cordic_CV.scala 67:42]
  wire [63:0] _current_theta_13_T_5 = $signed(current_theta_12) + 64'sh1ca5dc2; // @[Cordic_CV.scala 68:50]
  wire [49:0] _current_x_14_T = current_y_13[63:14]; // @[Cordic_CV.scala 62:62]
  wire [63:0] _GEN_97 = {{14{_current_x_14_T[49]}},_current_x_14_T}; // @[Cordic_CV.scala 62:42]
  wire [63:0] _current_x_14_T_3 = $signed(current_x_13) - $signed(_GEN_97); // @[Cordic_CV.scala 62:42]
  wire [63:0] _current_theta_14_T_2 = $signed(current_theta_13) - 64'she52ee1; // @[Cordic_CV.scala 64:50]
  wire [63:0] _current_x_14_T_7 = $signed(current_x_13) + $signed(_GEN_97); // @[Cordic_CV.scala 66:42]
  wire [63:0] _current_theta_14_T_5 = $signed(current_theta_13) + 64'she52ee1; // @[Cordic_CV.scala 68:50]
  wire [127:0] _io_r_T = $signed(current_x_14) * 64'sh9b74eda8; // @[Cordic_CV.scala 79:41]
  wire [95:0] _GEN_101 = _io_r_T[127:32]; // @[Cordic_CV.scala 79:8]
  assign io_theta = current_theta_14; // @[Cordic_CV.scala 78:12]
  assign io_r = _GEN_101[63:0]; // @[Cordic_CV.scala 79:8]
  always @(posedge clock) begin
    if (reset) begin // @[Cordic_CV.scala 40:43]
      current_x_0 <= 64'sh0; // @[Cordic_CV.scala 40:43]
    end else if ($signed(io_y) < 64'sh0) begin // @[Cordic_CV.scala 51:76]
      current_x_0 <= _current_x_0_T_3; // @[Cordic_CV.scala 52:22]
    end else begin
      current_x_0 <= _current_x_0_T_7; // @[Cordic_CV.scala 56:22]
    end
    if (reset) begin // @[Cordic_CV.scala 40:43]
      current_x_1 <= 64'sh0; // @[Cordic_CV.scala 40:43]
    end else if ($signed(current_y_0) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_x_1 <= _current_x_1_T_3; // @[Cordic_CV.scala 62:22]
    end else begin
      current_x_1 <= _current_x_1_T_7; // @[Cordic_CV.scala 66:22]
    end
    if (reset) begin // @[Cordic_CV.scala 40:43]
      current_x_2 <= 64'sh0; // @[Cordic_CV.scala 40:43]
    end else if ($signed(current_y_1) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_x_2 <= _current_x_2_T_3; // @[Cordic_CV.scala 62:22]
    end else begin
      current_x_2 <= _current_x_2_T_7; // @[Cordic_CV.scala 66:22]
    end
    if (reset) begin // @[Cordic_CV.scala 40:43]
      current_x_3 <= 64'sh0; // @[Cordic_CV.scala 40:43]
    end else if ($signed(current_y_2) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_x_3 <= _current_x_3_T_3; // @[Cordic_CV.scala 62:22]
    end else begin
      current_x_3 <= _current_x_3_T_7; // @[Cordic_CV.scala 66:22]
    end
    if (reset) begin // @[Cordic_CV.scala 40:43]
      current_x_4 <= 64'sh0; // @[Cordic_CV.scala 40:43]
    end else if ($signed(current_y_3) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_x_4 <= _current_x_4_T_3; // @[Cordic_CV.scala 62:22]
    end else begin
      current_x_4 <= _current_x_4_T_7; // @[Cordic_CV.scala 66:22]
    end
    if (reset) begin // @[Cordic_CV.scala 40:43]
      current_x_5 <= 64'sh0; // @[Cordic_CV.scala 40:43]
    end else if ($signed(current_y_4) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_x_5 <= _current_x_5_T_3; // @[Cordic_CV.scala 62:22]
    end else begin
      current_x_5 <= _current_x_5_T_7; // @[Cordic_CV.scala 66:22]
    end
    if (reset) begin // @[Cordic_CV.scala 40:43]
      current_x_6 <= 64'sh0; // @[Cordic_CV.scala 40:43]
    end else if ($signed(current_y_5) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_x_6 <= _current_x_6_T_3; // @[Cordic_CV.scala 62:22]
    end else begin
      current_x_6 <= _current_x_6_T_7; // @[Cordic_CV.scala 66:22]
    end
    if (reset) begin // @[Cordic_CV.scala 40:43]
      current_x_7 <= 64'sh0; // @[Cordic_CV.scala 40:43]
    end else if ($signed(current_y_6) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_x_7 <= _current_x_7_T_3; // @[Cordic_CV.scala 62:22]
    end else begin
      current_x_7 <= _current_x_7_T_7; // @[Cordic_CV.scala 66:22]
    end
    if (reset) begin // @[Cordic_CV.scala 40:43]
      current_x_8 <= 64'sh0; // @[Cordic_CV.scala 40:43]
    end else if ($signed(current_y_7) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_x_8 <= _current_x_8_T_3; // @[Cordic_CV.scala 62:22]
    end else begin
      current_x_8 <= _current_x_8_T_7; // @[Cordic_CV.scala 66:22]
    end
    if (reset) begin // @[Cordic_CV.scala 40:43]
      current_x_9 <= 64'sh0; // @[Cordic_CV.scala 40:43]
    end else if ($signed(current_y_8) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_x_9 <= _current_x_9_T_3; // @[Cordic_CV.scala 62:22]
    end else begin
      current_x_9 <= _current_x_9_T_7; // @[Cordic_CV.scala 66:22]
    end
    if (reset) begin // @[Cordic_CV.scala 40:43]
      current_x_10 <= 64'sh0; // @[Cordic_CV.scala 40:43]
    end else if ($signed(current_y_9) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_x_10 <= _current_x_10_T_3; // @[Cordic_CV.scala 62:22]
    end else begin
      current_x_10 <= _current_x_10_T_7; // @[Cordic_CV.scala 66:22]
    end
    if (reset) begin // @[Cordic_CV.scala 40:43]
      current_x_11 <= 64'sh0; // @[Cordic_CV.scala 40:43]
    end else if ($signed(current_y_10) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_x_11 <= _current_x_11_T_3; // @[Cordic_CV.scala 62:22]
    end else begin
      current_x_11 <= _current_x_11_T_7; // @[Cordic_CV.scala 66:22]
    end
    if (reset) begin // @[Cordic_CV.scala 40:43]
      current_x_12 <= 64'sh0; // @[Cordic_CV.scala 40:43]
    end else if ($signed(current_y_11) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_x_12 <= _current_x_12_T_3; // @[Cordic_CV.scala 62:22]
    end else begin
      current_x_12 <= _current_x_12_T_7; // @[Cordic_CV.scala 66:22]
    end
    if (reset) begin // @[Cordic_CV.scala 40:43]
      current_x_13 <= 64'sh0; // @[Cordic_CV.scala 40:43]
    end else if ($signed(current_y_12) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_x_13 <= _current_x_13_T_3; // @[Cordic_CV.scala 62:22]
    end else begin
      current_x_13 <= _current_x_13_T_7; // @[Cordic_CV.scala 66:22]
    end
    if (reset) begin // @[Cordic_CV.scala 40:43]
      current_x_14 <= 64'sh0; // @[Cordic_CV.scala 40:43]
    end else if ($signed(current_y_13) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_x_14 <= _current_x_14_T_3; // @[Cordic_CV.scala 62:22]
    end else begin
      current_x_14 <= _current_x_14_T_7; // @[Cordic_CV.scala 66:22]
    end
    if (reset) begin // @[Cordic_CV.scala 41:43]
      current_y_0 <= 64'sh0; // @[Cordic_CV.scala 41:43]
    end else if ($signed(io_y) < 64'sh0) begin // @[Cordic_CV.scala 51:76]
      current_y_0 <= _current_y_0_T_3; // @[Cordic_CV.scala 53:22]
    end else begin
      current_y_0 <= _current_y_0_T_7; // @[Cordic_CV.scala 57:22]
    end
    if (reset) begin // @[Cordic_CV.scala 41:43]
      current_y_1 <= 64'sh0; // @[Cordic_CV.scala 41:43]
    end else if ($signed(current_y_0) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_y_1 <= _current_y_1_T_3; // @[Cordic_CV.scala 63:22]
    end else begin
      current_y_1 <= _current_y_1_T_7; // @[Cordic_CV.scala 67:22]
    end
    if (reset) begin // @[Cordic_CV.scala 41:43]
      current_y_2 <= 64'sh0; // @[Cordic_CV.scala 41:43]
    end else if ($signed(current_y_1) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_y_2 <= _current_y_2_T_3; // @[Cordic_CV.scala 63:22]
    end else begin
      current_y_2 <= _current_y_2_T_7; // @[Cordic_CV.scala 67:22]
    end
    if (reset) begin // @[Cordic_CV.scala 41:43]
      current_y_3 <= 64'sh0; // @[Cordic_CV.scala 41:43]
    end else if ($signed(current_y_2) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_y_3 <= _current_y_3_T_3; // @[Cordic_CV.scala 63:22]
    end else begin
      current_y_3 <= _current_y_3_T_7; // @[Cordic_CV.scala 67:22]
    end
    if (reset) begin // @[Cordic_CV.scala 41:43]
      current_y_4 <= 64'sh0; // @[Cordic_CV.scala 41:43]
    end else if ($signed(current_y_3) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_y_4 <= _current_y_4_T_3; // @[Cordic_CV.scala 63:22]
    end else begin
      current_y_4 <= _current_y_4_T_7; // @[Cordic_CV.scala 67:22]
    end
    if (reset) begin // @[Cordic_CV.scala 41:43]
      current_y_5 <= 64'sh0; // @[Cordic_CV.scala 41:43]
    end else if ($signed(current_y_4) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_y_5 <= _current_y_5_T_3; // @[Cordic_CV.scala 63:22]
    end else begin
      current_y_5 <= _current_y_5_T_7; // @[Cordic_CV.scala 67:22]
    end
    if (reset) begin // @[Cordic_CV.scala 41:43]
      current_y_6 <= 64'sh0; // @[Cordic_CV.scala 41:43]
    end else if ($signed(current_y_5) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_y_6 <= _current_y_6_T_3; // @[Cordic_CV.scala 63:22]
    end else begin
      current_y_6 <= _current_y_6_T_7; // @[Cordic_CV.scala 67:22]
    end
    if (reset) begin // @[Cordic_CV.scala 41:43]
      current_y_7 <= 64'sh0; // @[Cordic_CV.scala 41:43]
    end else if ($signed(current_y_6) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_y_7 <= _current_y_7_T_3; // @[Cordic_CV.scala 63:22]
    end else begin
      current_y_7 <= _current_y_7_T_7; // @[Cordic_CV.scala 67:22]
    end
    if (reset) begin // @[Cordic_CV.scala 41:43]
      current_y_8 <= 64'sh0; // @[Cordic_CV.scala 41:43]
    end else if ($signed(current_y_7) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_y_8 <= _current_y_8_T_3; // @[Cordic_CV.scala 63:22]
    end else begin
      current_y_8 <= _current_y_8_T_7; // @[Cordic_CV.scala 67:22]
    end
    if (reset) begin // @[Cordic_CV.scala 41:43]
      current_y_9 <= 64'sh0; // @[Cordic_CV.scala 41:43]
    end else if ($signed(current_y_8) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_y_9 <= _current_y_9_T_3; // @[Cordic_CV.scala 63:22]
    end else begin
      current_y_9 <= _current_y_9_T_7; // @[Cordic_CV.scala 67:22]
    end
    if (reset) begin // @[Cordic_CV.scala 41:43]
      current_y_10 <= 64'sh0; // @[Cordic_CV.scala 41:43]
    end else if ($signed(current_y_9) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_y_10 <= _current_y_10_T_3; // @[Cordic_CV.scala 63:22]
    end else begin
      current_y_10 <= _current_y_10_T_7; // @[Cordic_CV.scala 67:22]
    end
    if (reset) begin // @[Cordic_CV.scala 41:43]
      current_y_11 <= 64'sh0; // @[Cordic_CV.scala 41:43]
    end else if ($signed(current_y_10) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_y_11 <= _current_y_11_T_3; // @[Cordic_CV.scala 63:22]
    end else begin
      current_y_11 <= _current_y_11_T_7; // @[Cordic_CV.scala 67:22]
    end
    if (reset) begin // @[Cordic_CV.scala 41:43]
      current_y_12 <= 64'sh0; // @[Cordic_CV.scala 41:43]
    end else if ($signed(current_y_11) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_y_12 <= _current_y_12_T_3; // @[Cordic_CV.scala 63:22]
    end else begin
      current_y_12 <= _current_y_12_T_7; // @[Cordic_CV.scala 67:22]
    end
    if (reset) begin // @[Cordic_CV.scala 41:43]
      current_y_13 <= 64'sh0; // @[Cordic_CV.scala 41:43]
    end else if ($signed(current_y_12) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_y_13 <= _current_y_13_T_3; // @[Cordic_CV.scala 63:22]
    end else begin
      current_y_13 <= _current_y_13_T_7; // @[Cordic_CV.scala 67:22]
    end
    if (reset) begin // @[Cordic_CV.scala 42:47]
      current_theta_0 <= 64'sh0; // @[Cordic_CV.scala 42:47]
    end else if ($signed(io_y) < 64'sh0) begin // @[Cordic_CV.scala 51:76]
      current_theta_0 <= _current_theta_0_T_2; // @[Cordic_CV.scala 54:26]
    end else begin
      current_theta_0 <= 64'sh2d00000000; // @[Cordic_CV.scala 58:26]
    end
    if (reset) begin // @[Cordic_CV.scala 42:47]
      current_theta_1 <= 64'sh0; // @[Cordic_CV.scala 42:47]
    end else if ($signed(current_y_0) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_theta_1 <= _current_theta_1_T_2; // @[Cordic_CV.scala 64:26]
    end else begin
      current_theta_1 <= _current_theta_1_T_5; // @[Cordic_CV.scala 68:26]
    end
    if (reset) begin // @[Cordic_CV.scala 42:47]
      current_theta_2 <= 64'sh0; // @[Cordic_CV.scala 42:47]
    end else if ($signed(current_y_1) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_theta_2 <= _current_theta_2_T_2; // @[Cordic_CV.scala 64:26]
    end else begin
      current_theta_2 <= _current_theta_2_T_5; // @[Cordic_CV.scala 68:26]
    end
    if (reset) begin // @[Cordic_CV.scala 42:47]
      current_theta_3 <= 64'sh0; // @[Cordic_CV.scala 42:47]
    end else if ($signed(current_y_2) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_theta_3 <= _current_theta_3_T_2; // @[Cordic_CV.scala 64:26]
    end else begin
      current_theta_3 <= _current_theta_3_T_5; // @[Cordic_CV.scala 68:26]
    end
    if (reset) begin // @[Cordic_CV.scala 42:47]
      current_theta_4 <= 64'sh0; // @[Cordic_CV.scala 42:47]
    end else if ($signed(current_y_3) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_theta_4 <= _current_theta_4_T_2; // @[Cordic_CV.scala 64:26]
    end else begin
      current_theta_4 <= _current_theta_4_T_5; // @[Cordic_CV.scala 68:26]
    end
    if (reset) begin // @[Cordic_CV.scala 42:47]
      current_theta_5 <= 64'sh0; // @[Cordic_CV.scala 42:47]
    end else if ($signed(current_y_4) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_theta_5 <= _current_theta_5_T_2; // @[Cordic_CV.scala 64:26]
    end else begin
      current_theta_5 <= _current_theta_5_T_5; // @[Cordic_CV.scala 68:26]
    end
    if (reset) begin // @[Cordic_CV.scala 42:47]
      current_theta_6 <= 64'sh0; // @[Cordic_CV.scala 42:47]
    end else if ($signed(current_y_5) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_theta_6 <= _current_theta_6_T_2; // @[Cordic_CV.scala 64:26]
    end else begin
      current_theta_6 <= _current_theta_6_T_5; // @[Cordic_CV.scala 68:26]
    end
    if (reset) begin // @[Cordic_CV.scala 42:47]
      current_theta_7 <= 64'sh0; // @[Cordic_CV.scala 42:47]
    end else if ($signed(current_y_6) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_theta_7 <= _current_theta_7_T_2; // @[Cordic_CV.scala 64:26]
    end else begin
      current_theta_7 <= _current_theta_7_T_5; // @[Cordic_CV.scala 68:26]
    end
    if (reset) begin // @[Cordic_CV.scala 42:47]
      current_theta_8 <= 64'sh0; // @[Cordic_CV.scala 42:47]
    end else if ($signed(current_y_7) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_theta_8 <= _current_theta_8_T_2; // @[Cordic_CV.scala 64:26]
    end else begin
      current_theta_8 <= _current_theta_8_T_5; // @[Cordic_CV.scala 68:26]
    end
    if (reset) begin // @[Cordic_CV.scala 42:47]
      current_theta_9 <= 64'sh0; // @[Cordic_CV.scala 42:47]
    end else if ($signed(current_y_8) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_theta_9 <= _current_theta_9_T_2; // @[Cordic_CV.scala 64:26]
    end else begin
      current_theta_9 <= _current_theta_9_T_5; // @[Cordic_CV.scala 68:26]
    end
    if (reset) begin // @[Cordic_CV.scala 42:47]
      current_theta_10 <= 64'sh0; // @[Cordic_CV.scala 42:47]
    end else if ($signed(current_y_9) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_theta_10 <= _current_theta_10_T_2; // @[Cordic_CV.scala 64:26]
    end else begin
      current_theta_10 <= _current_theta_10_T_5; // @[Cordic_CV.scala 68:26]
    end
    if (reset) begin // @[Cordic_CV.scala 42:47]
      current_theta_11 <= 64'sh0; // @[Cordic_CV.scala 42:47]
    end else if ($signed(current_y_10) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_theta_11 <= _current_theta_11_T_2; // @[Cordic_CV.scala 64:26]
    end else begin
      current_theta_11 <= _current_theta_11_T_5; // @[Cordic_CV.scala 68:26]
    end
    if (reset) begin // @[Cordic_CV.scala 42:47]
      current_theta_12 <= 64'sh0; // @[Cordic_CV.scala 42:47]
    end else if ($signed(current_y_11) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_theta_12 <= _current_theta_12_T_2; // @[Cordic_CV.scala 64:26]
    end else begin
      current_theta_12 <= _current_theta_12_T_5; // @[Cordic_CV.scala 68:26]
    end
    if (reset) begin // @[Cordic_CV.scala 42:47]
      current_theta_13 <= 64'sh0; // @[Cordic_CV.scala 42:47]
    end else if ($signed(current_y_12) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_theta_13 <= _current_theta_13_T_2; // @[Cordic_CV.scala 64:26]
    end else begin
      current_theta_13 <= _current_theta_13_T_5; // @[Cordic_CV.scala 68:26]
    end
    if (reset) begin // @[Cordic_CV.scala 42:47]
      current_theta_14 <= 64'sh0; // @[Cordic_CV.scala 42:47]
    end else if ($signed(current_y_13) < 64'sh0) begin // @[Cordic_CV.scala 61:88]
      current_theta_14 <= _current_theta_14_T_2; // @[Cordic_CV.scala 64:26]
    end else begin
      current_theta_14 <= _current_theta_14_T_5; // @[Cordic_CV.scala 68:26]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  current_x_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  current_x_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  current_x_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  current_x_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  current_x_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  current_x_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  current_x_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  current_x_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  current_x_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  current_x_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  current_x_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  current_x_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  current_x_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  current_x_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  current_x_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  current_y_0 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  current_y_1 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  current_y_2 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  current_y_3 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  current_y_4 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  current_y_5 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  current_y_6 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  current_y_7 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  current_y_8 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  current_y_9 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  current_y_10 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  current_y_11 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  current_y_12 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  current_y_13 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  current_theta_0 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  current_theta_1 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  current_theta_2 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  current_theta_3 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  current_theta_4 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  current_theta_5 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  current_theta_6 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  current_theta_7 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  current_theta_8 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  current_theta_9 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  current_theta_10 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  current_theta_11 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  current_theta_12 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  current_theta_13 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  current_theta_14 = _RAND_43[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cordic_cv(
  input         clock,
  input         reset,
  input  [63:0] io_x,
  input  [63:0] io_y,
  output [63:0] io_theta,
  output [63:0] io_r
);
  wire  cordic_cv_unit_clock; // @[Cordic_CV.scala 104:30]
  wire  cordic_cv_unit_reset; // @[Cordic_CV.scala 104:30]
  wire [63:0] cordic_cv_unit_io_x; // @[Cordic_CV.scala 104:30]
  wire [63:0] cordic_cv_unit_io_y; // @[Cordic_CV.scala 104:30]
  wire [63:0] cordic_cv_unit_io_theta; // @[Cordic_CV.scala 104:30]
  wire [63:0] cordic_cv_unit_io_r; // @[Cordic_CV.scala 104:30]
  wire [63:0] _cordic_cv_unit_io_x_T_2 = 64'sh0 - $signed(io_x); // @[Cordic_CV.scala 107:28]
  wire [63:0] _cordic_cv_unit_io_y_T_2 = 64'sh0 - $signed(io_y); // @[Cordic_CV.scala 108:28]
  wire [63:0] _io_theta_T_2 = $signed(cordic_cv_unit_io_theta) + 64'shb400000000; // @[Cordic_CV.scala 110:43]
  wire [63:0] _io_theta_T_5 = $signed(cordic_cv_unit_io_theta) - 64'shb400000000; // @[Cordic_CV.scala 112:43]
  wire [63:0] _GEN_0 = $signed(io_y) > 64'sh0 ? $signed(_io_theta_T_2) : $signed(_io_theta_T_5); // @[Cordic_CV.scala 109:71 110:16 112:16]
  CORDIC_CV_ORIGIN cordic_cv_unit ( // @[Cordic_CV.scala 104:30]
    .clock(cordic_cv_unit_clock),
    .reset(cordic_cv_unit_reset),
    .io_x(cordic_cv_unit_io_x),
    .io_y(cordic_cv_unit_io_y),
    .io_theta(cordic_cv_unit_io_theta),
    .io_r(cordic_cv_unit_io_r)
  );
  assign io_theta = $signed(io_x) < 64'sh0 ? $signed(_GEN_0) : $signed(cordic_cv_unit_io_theta); // @[Cordic_CV.scala 106:69 117:14]
  assign io_r = cordic_cv_unit_io_r; // @[Cordic_CV.scala 120:8]
  assign cordic_cv_unit_clock = clock;
  assign cordic_cv_unit_reset = reset;
  assign cordic_cv_unit_io_x = $signed(io_x) < 64'sh0 ? $signed(_cordic_cv_unit_io_x_T_2) : $signed(io_x); // @[Cordic_CV.scala 106:69 107:25 115:25]
  assign cordic_cv_unit_io_y = $signed(io_x) < 64'sh0 ? $signed(_cordic_cv_unit_io_y_T_2) : $signed(io_y); // @[Cordic_CV.scala 106:69 108:25 116:25]
endmodule
module cordic_complex_divide(
  input         clock,
  input         reset,
  input  [63:0] io_op2_re,
  input  [63:0] io_op2_im,
  output [63:0] io_res_re,
  output [63:0] io_res_im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
`endif // RANDOMIZE_REG_INIT
  wire  cordic_cv_clock; // @[Cordic_CV.scala 141:27]
  wire  cordic_cv_reset; // @[Cordic_CV.scala 141:27]
  wire [63:0] cordic_cv_io_x; // @[Cordic_CV.scala 141:27]
  wire [63:0] cordic_cv_io_y; // @[Cordic_CV.scala 141:27]
  wire [63:0] cordic_cv_io_theta; // @[Cordic_CV.scala 141:27]
  wire [63:0] cordic_cv_io_r; // @[Cordic_CV.scala 141:27]
  wire  z_a_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  z_a_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] z_a_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] z_a_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] z_a_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  z_b_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  z_b_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] z_b_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] z_b_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] z_b_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  cordic_unit_clock; // @[Cordic_CR.scala 96:47]
  wire  cordic_unit_reset; // @[Cordic_CR.scala 96:47]
  wire [63:0] cordic_unit_io_x; // @[Cordic_CR.scala 96:47]
  wire [63:0] cordic_unit_io_y; // @[Cordic_CR.scala 96:47]
  wire [63:0] cordic_unit_io_theta; // @[Cordic_CR.scala 96:47]
  wire [63:0] cordic_unit_io_x_n; // @[Cordic_CR.scala 96:47]
  wire [63:0] cordic_unit_io_y_n; // @[Cordic_CR.scala 96:47]
  reg  flag_reg_0; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_1; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_2; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_3; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_4; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_5; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_6; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_7; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_8; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_9; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_10; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_11; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_12; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_13; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_14; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_15; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_16; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_17; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_18; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_19; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_20; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_21; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_22; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_23; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_24; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_25; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_26; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_27; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_28; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_29; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_30; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_31; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_32; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_33; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_34; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_35; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_36; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_37; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_38; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_39; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_40; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_41; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_42; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_43; // @[Cordic_Complex_Divide.scala 19:36]
  reg  flag_reg_44; // @[Cordic_Complex_Divide.scala 19:36]
  wire [63:0] _p_T_2 = 64'sh0 - $signed(io_op2_re); // @[Cordic_Complex_Divide.scala 21:10]
  wire [63:0] _q_T_2 = 64'sh0 - $signed(io_op2_im); // @[Cordic_Complex_Divide.scala 22:10]
  wire  _GEN_2 = $signed(io_op2_re) < 64'sh0 ? 1'h0 : 1'h1; // @[Cordic_Complex_Divide.scala 20:75 23:17 27:17]
  reg [63:0] a_reg_0; // @[Cordic_Complex_Divide.scala 34:39]
  reg [63:0] a_reg_1; // @[Cordic_Complex_Divide.scala 34:39]
  reg [63:0] a_reg_2; // @[Cordic_Complex_Divide.scala 34:39]
  reg [63:0] a_reg_3; // @[Cordic_Complex_Divide.scala 34:39]
  reg [63:0] a_reg_4; // @[Cordic_Complex_Divide.scala 34:39]
  reg [63:0] a_reg_5; // @[Cordic_Complex_Divide.scala 34:39]
  reg [63:0] a_reg_6; // @[Cordic_Complex_Divide.scala 34:39]
  reg [63:0] a_reg_7; // @[Cordic_Complex_Divide.scala 34:39]
  reg [63:0] a_reg_8; // @[Cordic_Complex_Divide.scala 34:39]
  reg [63:0] a_reg_9; // @[Cordic_Complex_Divide.scala 34:39]
  reg [63:0] a_reg_10; // @[Cordic_Complex_Divide.scala 34:39]
  reg [63:0] a_reg_11; // @[Cordic_Complex_Divide.scala 34:39]
  reg [63:0] a_reg_12; // @[Cordic_Complex_Divide.scala 34:39]
  reg [63:0] a_reg_13; // @[Cordic_Complex_Divide.scala 34:39]
  reg [63:0] a_reg_14; // @[Cordic_Complex_Divide.scala 34:39]
  reg [63:0] theta_reg_0; // @[Cordic_Complex_Divide.scala 50:43]
  reg [63:0] theta_reg_1; // @[Cordic_Complex_Divide.scala 50:43]
  reg [63:0] theta_reg_2; // @[Cordic_Complex_Divide.scala 50:43]
  reg [63:0] theta_reg_3; // @[Cordic_Complex_Divide.scala 50:43]
  reg [63:0] theta_reg_4; // @[Cordic_Complex_Divide.scala 50:43]
  reg [63:0] theta_reg_5; // @[Cordic_Complex_Divide.scala 50:43]
  reg [63:0] theta_reg_6; // @[Cordic_Complex_Divide.scala 50:43]
  reg [63:0] theta_reg_7; // @[Cordic_Complex_Divide.scala 50:43]
  reg [63:0] theta_reg_8; // @[Cordic_Complex_Divide.scala 50:43]
  reg [63:0] theta_reg_9; // @[Cordic_Complex_Divide.scala 50:43]
  reg [63:0] theta_reg_10; // @[Cordic_Complex_Divide.scala 50:43]
  reg [63:0] theta_reg_11; // @[Cordic_Complex_Divide.scala 50:43]
  reg [63:0] theta_reg_12; // @[Cordic_Complex_Divide.scala 50:43]
  reg [63:0] theta_reg_13; // @[Cordic_Complex_Divide.scala 50:43]
  reg [63:0] theta_reg_14; // @[Cordic_Complex_Divide.scala 50:43]
  wire [63:0] _io_res_re_T_2 = 64'sh0 - $signed(cordic_unit_io_x_n); // @[Cordic_Complex_Divide.scala 70:18]
  wire [63:0] _io_res_im_T_2 = 64'sh0 - $signed(cordic_unit_io_y_n); // @[Cordic_Complex_Divide.scala 71:18]
  cordic_cv cordic_cv ( // @[Cordic_CV.scala 141:27]
    .clock(cordic_cv_clock),
    .reset(cordic_cv_reset),
    .io_x(cordic_cv_io_x),
    .io_y(cordic_cv_io_y),
    .io_theta(cordic_cv_io_theta),
    .io_r(cordic_cv_io_r)
  );
  cordic_divide z_a_divide ( // @[Cordic_LV.scala 211:24]
    .clock(z_a_divide_clock),
    .reset(z_a_divide_reset),
    .io_x(z_a_divide_io_x),
    .io_y(z_a_divide_io_y),
    .io_z(z_a_divide_io_z)
  );
  cordic_divide z_b_divide ( // @[Cordic_LV.scala 211:24]
    .clock(z_b_divide_clock),
    .reset(z_b_divide_reset),
    .io_x(z_b_divide_io_x),
    .io_y(z_b_divide_io_y),
    .io_z(z_b_divide_io_z)
  );
  CORDIC_CR_ORIGIN cordic_unit ( // @[Cordic_CR.scala 96:47]
    .clock(cordic_unit_clock),
    .reset(cordic_unit_reset),
    .io_x(cordic_unit_io_x),
    .io_y(cordic_unit_io_y),
    .io_theta(cordic_unit_io_theta),
    .io_x_n(cordic_unit_io_x_n),
    .io_y_n(cordic_unit_io_y_n)
  );
  assign io_res_re = flag_reg_44 ? $signed(cordic_unit_io_x_n) : $signed(_io_res_re_T_2); // @[Cordic_Complex_Divide.scala 66:42 67:15 70:15]
  assign io_res_im = flag_reg_44 ? $signed(cordic_unit_io_y_n) : $signed(_io_res_im_T_2); // @[Cordic_Complex_Divide.scala 66:42 68:15 71:15]
  assign cordic_cv_clock = clock;
  assign cordic_cv_reset = reset;
  assign cordic_cv_io_x = $signed(io_op2_re) < 64'sh0 ? $signed(_p_T_2) : $signed(io_op2_re); // @[Cordic_Complex_Divide.scala 20:75 21:7 25:7]
  assign cordic_cv_io_y = $signed(io_op2_re) < 64'sh0 ? $signed(_q_T_2) : $signed(io_op2_im); // @[Cordic_Complex_Divide.scala 20:75 22:7 26:7]
  assign z_a_divide_clock = clock;
  assign z_a_divide_reset = reset;
  assign z_a_divide_io_x = cordic_cv_io_r; // @[Cordic_LV.scala 212:17]
  assign z_a_divide_io_y = a_reg_14; // @[Cordic_LV.scala 213:17]
  assign z_b_divide_clock = clock;
  assign z_b_divide_reset = reset;
  assign z_b_divide_io_x = cordic_cv_io_r; // @[Cordic_LV.scala 212:17]
  assign z_b_divide_io_y = 64'sh0; // @[Cordic_LV.scala 213:17]
  assign cordic_unit_clock = clock;
  assign cordic_unit_reset = reset;
  assign cordic_unit_io_x = z_a_divide_io_z; // @[Cordic_CR.scala 97:22]
  assign cordic_unit_io_y = z_b_divide_io_z; // @[Cordic_CR.scala 98:22]
  assign cordic_unit_io_theta = 64'sh0 - $signed(theta_reg_14); // @[Cordic_Complex_Divide.scala 64:38]
  always @(posedge clock) begin
    flag_reg_0 <= reset | _GEN_2; // @[Cordic_Complex_Divide.scala 19:{36,36}]
    flag_reg_1 <= reset | flag_reg_0; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_2 <= reset | flag_reg_1; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_3 <= reset | flag_reg_2; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_4 <= reset | flag_reg_3; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_5 <= reset | flag_reg_4; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_6 <= reset | flag_reg_5; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_7 <= reset | flag_reg_6; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_8 <= reset | flag_reg_7; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_9 <= reset | flag_reg_8; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_10 <= reset | flag_reg_9; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_11 <= reset | flag_reg_10; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_12 <= reset | flag_reg_11; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_13 <= reset | flag_reg_12; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_14 <= reset | flag_reg_13; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_15 <= reset | flag_reg_14; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_16 <= reset | flag_reg_15; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_17 <= reset | flag_reg_16; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_18 <= reset | flag_reg_17; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_19 <= reset | flag_reg_18; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_20 <= reset | flag_reg_19; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_21 <= reset | flag_reg_20; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_22 <= reset | flag_reg_21; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_23 <= reset | flag_reg_22; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_24 <= reset | flag_reg_23; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_25 <= reset | flag_reg_24; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_26 <= reset | flag_reg_25; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_27 <= reset | flag_reg_26; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_28 <= reset | flag_reg_27; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_29 <= reset | flag_reg_28; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_30 <= reset | flag_reg_29; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_31 <= reset | flag_reg_30; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_32 <= reset | flag_reg_31; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_33 <= reset | flag_reg_32; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_34 <= reset | flag_reg_33; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_35 <= reset | flag_reg_34; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_36 <= reset | flag_reg_35; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_37 <= reset | flag_reg_36; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_38 <= reset | flag_reg_37; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_39 <= reset | flag_reg_38; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_40 <= reset | flag_reg_39; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_41 <= reset | flag_reg_40; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_42 <= reset | flag_reg_41; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_43 <= reset | flag_reg_42; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    flag_reg_44 <= reset | flag_reg_43; // @[Cordic_Complex_Divide.scala 19:{36,36} 30:17]
    if (reset) begin // @[Cordic_Complex_Divide.scala 34:39]
      a_reg_0 <= 64'sh0; // @[Cordic_Complex_Divide.scala 34:39]
    end else begin
      a_reg_0 <= 64'sh100000000; // @[Cordic_Complex_Divide.scala 38:16]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 34:39]
      a_reg_1 <= 64'sh0; // @[Cordic_Complex_Divide.scala 34:39]
    end else begin
      a_reg_1 <= a_reg_0; // @[Cordic_Complex_Divide.scala 41:16]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 34:39]
      a_reg_2 <= 64'sh0; // @[Cordic_Complex_Divide.scala 34:39]
    end else begin
      a_reg_2 <= a_reg_1; // @[Cordic_Complex_Divide.scala 41:16]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 34:39]
      a_reg_3 <= 64'sh0; // @[Cordic_Complex_Divide.scala 34:39]
    end else begin
      a_reg_3 <= a_reg_2; // @[Cordic_Complex_Divide.scala 41:16]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 34:39]
      a_reg_4 <= 64'sh0; // @[Cordic_Complex_Divide.scala 34:39]
    end else begin
      a_reg_4 <= a_reg_3; // @[Cordic_Complex_Divide.scala 41:16]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 34:39]
      a_reg_5 <= 64'sh0; // @[Cordic_Complex_Divide.scala 34:39]
    end else begin
      a_reg_5 <= a_reg_4; // @[Cordic_Complex_Divide.scala 41:16]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 34:39]
      a_reg_6 <= 64'sh0; // @[Cordic_Complex_Divide.scala 34:39]
    end else begin
      a_reg_6 <= a_reg_5; // @[Cordic_Complex_Divide.scala 41:16]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 34:39]
      a_reg_7 <= 64'sh0; // @[Cordic_Complex_Divide.scala 34:39]
    end else begin
      a_reg_7 <= a_reg_6; // @[Cordic_Complex_Divide.scala 41:16]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 34:39]
      a_reg_8 <= 64'sh0; // @[Cordic_Complex_Divide.scala 34:39]
    end else begin
      a_reg_8 <= a_reg_7; // @[Cordic_Complex_Divide.scala 41:16]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 34:39]
      a_reg_9 <= 64'sh0; // @[Cordic_Complex_Divide.scala 34:39]
    end else begin
      a_reg_9 <= a_reg_8; // @[Cordic_Complex_Divide.scala 41:16]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 34:39]
      a_reg_10 <= 64'sh0; // @[Cordic_Complex_Divide.scala 34:39]
    end else begin
      a_reg_10 <= a_reg_9; // @[Cordic_Complex_Divide.scala 41:16]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 34:39]
      a_reg_11 <= 64'sh0; // @[Cordic_Complex_Divide.scala 34:39]
    end else begin
      a_reg_11 <= a_reg_10; // @[Cordic_Complex_Divide.scala 41:16]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 34:39]
      a_reg_12 <= 64'sh0; // @[Cordic_Complex_Divide.scala 34:39]
    end else begin
      a_reg_12 <= a_reg_11; // @[Cordic_Complex_Divide.scala 41:16]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 34:39]
      a_reg_13 <= 64'sh0; // @[Cordic_Complex_Divide.scala 34:39]
    end else begin
      a_reg_13 <= a_reg_12; // @[Cordic_Complex_Divide.scala 41:16]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 34:39]
      a_reg_14 <= 64'sh0; // @[Cordic_Complex_Divide.scala 34:39]
    end else begin
      a_reg_14 <= a_reg_13; // @[Cordic_Complex_Divide.scala 41:16]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 50:43]
      theta_reg_0 <= 64'sh0; // @[Cordic_Complex_Divide.scala 50:43]
    end else begin
      theta_reg_0 <= cordic_cv_io_theta; // @[Cordic_Complex_Divide.scala 53:20]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 50:43]
      theta_reg_1 <= 64'sh0; // @[Cordic_Complex_Divide.scala 50:43]
    end else begin
      theta_reg_1 <= theta_reg_0; // @[Cordic_Complex_Divide.scala 55:20]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 50:43]
      theta_reg_2 <= 64'sh0; // @[Cordic_Complex_Divide.scala 50:43]
    end else begin
      theta_reg_2 <= theta_reg_1; // @[Cordic_Complex_Divide.scala 55:20]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 50:43]
      theta_reg_3 <= 64'sh0; // @[Cordic_Complex_Divide.scala 50:43]
    end else begin
      theta_reg_3 <= theta_reg_2; // @[Cordic_Complex_Divide.scala 55:20]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 50:43]
      theta_reg_4 <= 64'sh0; // @[Cordic_Complex_Divide.scala 50:43]
    end else begin
      theta_reg_4 <= theta_reg_3; // @[Cordic_Complex_Divide.scala 55:20]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 50:43]
      theta_reg_5 <= 64'sh0; // @[Cordic_Complex_Divide.scala 50:43]
    end else begin
      theta_reg_5 <= theta_reg_4; // @[Cordic_Complex_Divide.scala 55:20]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 50:43]
      theta_reg_6 <= 64'sh0; // @[Cordic_Complex_Divide.scala 50:43]
    end else begin
      theta_reg_6 <= theta_reg_5; // @[Cordic_Complex_Divide.scala 55:20]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 50:43]
      theta_reg_7 <= 64'sh0; // @[Cordic_Complex_Divide.scala 50:43]
    end else begin
      theta_reg_7 <= theta_reg_6; // @[Cordic_Complex_Divide.scala 55:20]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 50:43]
      theta_reg_8 <= 64'sh0; // @[Cordic_Complex_Divide.scala 50:43]
    end else begin
      theta_reg_8 <= theta_reg_7; // @[Cordic_Complex_Divide.scala 55:20]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 50:43]
      theta_reg_9 <= 64'sh0; // @[Cordic_Complex_Divide.scala 50:43]
    end else begin
      theta_reg_9 <= theta_reg_8; // @[Cordic_Complex_Divide.scala 55:20]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 50:43]
      theta_reg_10 <= 64'sh0; // @[Cordic_Complex_Divide.scala 50:43]
    end else begin
      theta_reg_10 <= theta_reg_9; // @[Cordic_Complex_Divide.scala 55:20]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 50:43]
      theta_reg_11 <= 64'sh0; // @[Cordic_Complex_Divide.scala 50:43]
    end else begin
      theta_reg_11 <= theta_reg_10; // @[Cordic_Complex_Divide.scala 55:20]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 50:43]
      theta_reg_12 <= 64'sh0; // @[Cordic_Complex_Divide.scala 50:43]
    end else begin
      theta_reg_12 <= theta_reg_11; // @[Cordic_Complex_Divide.scala 55:20]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 50:43]
      theta_reg_13 <= 64'sh0; // @[Cordic_Complex_Divide.scala 50:43]
    end else begin
      theta_reg_13 <= theta_reg_12; // @[Cordic_Complex_Divide.scala 55:20]
    end
    if (reset) begin // @[Cordic_Complex_Divide.scala 50:43]
      theta_reg_14 <= 64'sh0; // @[Cordic_Complex_Divide.scala 50:43]
    end else begin
      theta_reg_14 <= theta_reg_13; // @[Cordic_Complex_Divide.scala 55:20]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flag_reg_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  flag_reg_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  flag_reg_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  flag_reg_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  flag_reg_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  flag_reg_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  flag_reg_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  flag_reg_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  flag_reg_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  flag_reg_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  flag_reg_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  flag_reg_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  flag_reg_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  flag_reg_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  flag_reg_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  flag_reg_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  flag_reg_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  flag_reg_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  flag_reg_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  flag_reg_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  flag_reg_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  flag_reg_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  flag_reg_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  flag_reg_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  flag_reg_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  flag_reg_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  flag_reg_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  flag_reg_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  flag_reg_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  flag_reg_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  flag_reg_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  flag_reg_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  flag_reg_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  flag_reg_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  flag_reg_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  flag_reg_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  flag_reg_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  flag_reg_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  flag_reg_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  flag_reg_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  flag_reg_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  flag_reg_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  flag_reg_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  flag_reg_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  flag_reg_44 = _RAND_44[0:0];
  _RAND_45 = {2{`RANDOM}};
  a_reg_0 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  a_reg_1 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  a_reg_2 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  a_reg_3 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  a_reg_4 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  a_reg_5 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  a_reg_6 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  a_reg_7 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  a_reg_8 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  a_reg_9 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  a_reg_10 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  a_reg_11 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  a_reg_12 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  a_reg_13 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  a_reg_14 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  theta_reg_0 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  theta_reg_1 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  theta_reg_2 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  theta_reg_3 = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  theta_reg_4 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  theta_reg_5 = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  theta_reg_6 = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  theta_reg_7 = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  theta_reg_8 = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  theta_reg_9 = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  theta_reg_10 = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  theta_reg_11 = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  theta_reg_12 = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  theta_reg_13 = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  theta_reg_14 = _RAND_74[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module matrix_mul_v1_1(
  input         clock,
  input         io_reset,
  input         io_ready,
  input  [63:0] io_matrixA_0_re,
  input  [63:0] io_matrixA_0_im,
  input  [63:0] io_matrixA_1_re,
  input  [63:0] io_matrixA_1_im,
  input  [63:0] io_matrixA_2_re,
  input  [63:0] io_matrixA_2_im,
  input  [63:0] io_matrixB_0_re,
  input  [63:0] io_matrixB_0_im,
  input  [63:0] io_matrixB_1_re,
  input  [63:0] io_matrixB_1_im,
  input  [63:0] io_matrixB_2_re,
  input  [63:0] io_matrixB_2_im,
  output [63:0] io_matrixC_0_re,
  output [63:0] io_matrixC_0_im,
  output [63:0] io_matrixC_1_re,
  output [63:0] io_matrixC_1_im,
  output [63:0] io_matrixC_2_re,
  output [63:0] io_matrixC_2_im,
  output [63:0] io_matrixC_3_re,
  output [63:0] io_matrixC_3_im,
  output [63:0] io_matrixC_4_re,
  output [63:0] io_matrixC_4_im,
  output [63:0] io_matrixC_5_re,
  output [63:0] io_matrixC_5_im,
  output [63:0] io_matrixC_6_re,
  output [63:0] io_matrixC_6_im,
  output [63:0] io_matrixC_7_re,
  output [63:0] io_matrixC_7_im,
  output [63:0] io_matrixC_8_re,
  output [63:0] io_matrixC_8_im,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  PE_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_1_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_1_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_2_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_2_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_3_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_3_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_4_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_4_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_5_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_5_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_6_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_6_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_7_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_7_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_8_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_8_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  reg [63:0] regsA_0_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_0_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_1_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_1_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_2_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_2_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsB_0_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_0_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_1_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_1_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_2_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_2_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [3:0] input_point; // @[Matrix_Mul_V1.scala 84:30]
  wire [3:0] _input_point_T_1 = input_point + 4'h1; // @[Matrix_Mul_V1.scala 116:32]
  wire  _T = input_point < 4'h3; // @[Matrix_Mul_V1.scala 145:20]
  wire [2:0] _T_1 = 1'h0 * 2'h3; // @[Matrix_Mul_V1.scala 148:44]
  wire [3:0] _GEN_149 = {{1'd0}, _T_1}; // @[Matrix_Mul_V1.scala 148:60]
  wire [3:0] _T_3 = _GEN_149 + input_point; // @[Matrix_Mul_V1.scala 148:60]
  wire [63:0] _GEN_29 = 4'h1 == _T_3 ? $signed(64'sh0) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_30 = 4'h2 == _T_3 ? $signed(64'sh0) : $signed(_GEN_29); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_31 = 4'h3 == _T_3 ? $signed(64'sh0) : $signed(_GEN_30); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_32 = 4'h4 == _T_3 ? $signed(regsA_1_im) : $signed(_GEN_31); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_33 = 4'h5 == _T_3 ? $signed(64'sh0) : $signed(_GEN_32); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_34 = 4'h6 == _T_3 ? $signed(64'sh0) : $signed(_GEN_33); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_35 = 4'h7 == _T_3 ? $signed(64'sh0) : $signed(_GEN_34); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_36 = 4'h8 == _T_3 ? $signed(regsA_2_im) : $signed(_GEN_35); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_38 = 4'h1 == _T_3 ? $signed(64'sh0) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_39 = 4'h2 == _T_3 ? $signed(64'sh0) : $signed(_GEN_38); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_40 = 4'h3 == _T_3 ? $signed(64'sh0) : $signed(_GEN_39); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_41 = 4'h4 == _T_3 ? $signed(regsA_1_re) : $signed(_GEN_40); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_42 = 4'h5 == _T_3 ? $signed(64'sh0) : $signed(_GEN_41); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_43 = 4'h6 == _T_3 ? $signed(64'sh0) : $signed(_GEN_42); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_44 = 4'h7 == _T_3 ? $signed(64'sh0) : $signed(_GEN_43); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_45 = 4'h8 == _T_3 ? $signed(regsA_2_re) : $signed(_GEN_44); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [2:0] _T_4 = 1'h1 * 2'h3; // @[Matrix_Mul_V1.scala 148:44]
  wire [3:0] _GEN_150 = {{1'd0}, _T_4}; // @[Matrix_Mul_V1.scala 148:60]
  wire [3:0] _T_6 = _GEN_150 + input_point; // @[Matrix_Mul_V1.scala 148:60]
  wire [63:0] _GEN_47 = 4'h1 == _T_6 ? $signed(64'sh0) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_48 = 4'h2 == _T_6 ? $signed(64'sh0) : $signed(_GEN_47); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_49 = 4'h3 == _T_6 ? $signed(64'sh0) : $signed(_GEN_48); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_50 = 4'h4 == _T_6 ? $signed(regsA_1_im) : $signed(_GEN_49); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_51 = 4'h5 == _T_6 ? $signed(64'sh0) : $signed(_GEN_50); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_52 = 4'h6 == _T_6 ? $signed(64'sh0) : $signed(_GEN_51); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_53 = 4'h7 == _T_6 ? $signed(64'sh0) : $signed(_GEN_52); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_54 = 4'h8 == _T_6 ? $signed(regsA_2_im) : $signed(_GEN_53); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_56 = 4'h1 == _T_6 ? $signed(64'sh0) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_57 = 4'h2 == _T_6 ? $signed(64'sh0) : $signed(_GEN_56); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_58 = 4'h3 == _T_6 ? $signed(64'sh0) : $signed(_GEN_57); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_59 = 4'h4 == _T_6 ? $signed(regsA_1_re) : $signed(_GEN_58); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_60 = 4'h5 == _T_6 ? $signed(64'sh0) : $signed(_GEN_59); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_61 = 4'h6 == _T_6 ? $signed(64'sh0) : $signed(_GEN_60); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_62 = 4'h7 == _T_6 ? $signed(64'sh0) : $signed(_GEN_61); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_63 = 4'h8 == _T_6 ? $signed(regsA_2_re) : $signed(_GEN_62); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [3:0] _T_7 = 2'h2 * 2'h3; // @[Matrix_Mul_V1.scala 148:44]
  wire [3:0] _T_9 = _T_7 + input_point; // @[Matrix_Mul_V1.scala 148:60]
  wire [63:0] _GEN_65 = 4'h1 == _T_9 ? $signed(64'sh0) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_66 = 4'h2 == _T_9 ? $signed(64'sh0) : $signed(_GEN_65); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_67 = 4'h3 == _T_9 ? $signed(64'sh0) : $signed(_GEN_66); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_68 = 4'h4 == _T_9 ? $signed(regsA_1_im) : $signed(_GEN_67); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_69 = 4'h5 == _T_9 ? $signed(64'sh0) : $signed(_GEN_68); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_70 = 4'h6 == _T_9 ? $signed(64'sh0) : $signed(_GEN_69); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_71 = 4'h7 == _T_9 ? $signed(64'sh0) : $signed(_GEN_70); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_72 = 4'h8 == _T_9 ? $signed(regsA_2_im) : $signed(_GEN_71); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_74 = 4'h1 == _T_9 ? $signed(64'sh0) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_75 = 4'h2 == _T_9 ? $signed(64'sh0) : $signed(_GEN_74); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_76 = 4'h3 == _T_9 ? $signed(64'sh0) : $signed(_GEN_75); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_77 = 4'h4 == _T_9 ? $signed(regsA_1_re) : $signed(_GEN_76); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_78 = 4'h5 == _T_9 ? $signed(64'sh0) : $signed(_GEN_77); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_79 = 4'h6 == _T_9 ? $signed(64'sh0) : $signed(_GEN_78); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_80 = 4'h7 == _T_9 ? $signed(64'sh0) : $signed(_GEN_79); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_81 = 4'h8 == _T_9 ? $signed(regsA_2_re) : $signed(_GEN_80); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_89 = 4'h1 == _T_3 ? $signed(64'sh0) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_90 = 4'h2 == _T_3 ? $signed(64'sh0) : $signed(_GEN_89); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_91 = 4'h3 == _T_3 ? $signed(64'sh0) : $signed(_GEN_90); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_92 = 4'h4 == _T_3 ? $signed(regsB_1_im) : $signed(_GEN_91); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_93 = 4'h5 == _T_3 ? $signed(64'sh0) : $signed(_GEN_92); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_94 = 4'h6 == _T_3 ? $signed(64'sh0) : $signed(_GEN_93); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_95 = 4'h7 == _T_3 ? $signed(64'sh0) : $signed(_GEN_94); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_96 = 4'h8 == _T_3 ? $signed(regsB_2_im) : $signed(_GEN_95); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_98 = 4'h1 == _T_3 ? $signed(64'sh0) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_99 = 4'h2 == _T_3 ? $signed(64'sh0) : $signed(_GEN_98); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_100 = 4'h3 == _T_3 ? $signed(64'sh0) : $signed(_GEN_99); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_101 = 4'h4 == _T_3 ? $signed(regsB_1_re) : $signed(_GEN_100); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_102 = 4'h5 == _T_3 ? $signed(64'sh0) : $signed(_GEN_101); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_103 = 4'h6 == _T_3 ? $signed(64'sh0) : $signed(_GEN_102); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_104 = 4'h7 == _T_3 ? $signed(64'sh0) : $signed(_GEN_103); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_105 = 4'h8 == _T_3 ? $signed(regsB_2_re) : $signed(_GEN_104); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_107 = 4'h1 == _T_6 ? $signed(64'sh0) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_108 = 4'h2 == _T_6 ? $signed(64'sh0) : $signed(_GEN_107); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_109 = 4'h3 == _T_6 ? $signed(64'sh0) : $signed(_GEN_108); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_110 = 4'h4 == _T_6 ? $signed(regsB_1_im) : $signed(_GEN_109); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_111 = 4'h5 == _T_6 ? $signed(64'sh0) : $signed(_GEN_110); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_112 = 4'h6 == _T_6 ? $signed(64'sh0) : $signed(_GEN_111); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_113 = 4'h7 == _T_6 ? $signed(64'sh0) : $signed(_GEN_112); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_114 = 4'h8 == _T_6 ? $signed(regsB_2_im) : $signed(_GEN_113); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_116 = 4'h1 == _T_6 ? $signed(64'sh0) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_117 = 4'h2 == _T_6 ? $signed(64'sh0) : $signed(_GEN_116); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_118 = 4'h3 == _T_6 ? $signed(64'sh0) : $signed(_GEN_117); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_119 = 4'h4 == _T_6 ? $signed(regsB_1_re) : $signed(_GEN_118); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_120 = 4'h5 == _T_6 ? $signed(64'sh0) : $signed(_GEN_119); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_121 = 4'h6 == _T_6 ? $signed(64'sh0) : $signed(_GEN_120); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_122 = 4'h7 == _T_6 ? $signed(64'sh0) : $signed(_GEN_121); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_123 = 4'h8 == _T_6 ? $signed(regsB_2_re) : $signed(_GEN_122); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_125 = 4'h1 == _T_9 ? $signed(64'sh0) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_126 = 4'h2 == _T_9 ? $signed(64'sh0) : $signed(_GEN_125); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_127 = 4'h3 == _T_9 ? $signed(64'sh0) : $signed(_GEN_126); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_128 = 4'h4 == _T_9 ? $signed(regsB_1_im) : $signed(_GEN_127); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_129 = 4'h5 == _T_9 ? $signed(64'sh0) : $signed(_GEN_128); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_130 = 4'h6 == _T_9 ? $signed(64'sh0) : $signed(_GEN_129); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_131 = 4'h7 == _T_9 ? $signed(64'sh0) : $signed(_GEN_130); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_132 = 4'h8 == _T_9 ? $signed(regsB_2_im) : $signed(_GEN_131); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_134 = 4'h1 == _T_9 ? $signed(64'sh0) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_135 = 4'h2 == _T_9 ? $signed(64'sh0) : $signed(_GEN_134); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_136 = 4'h3 == _T_9 ? $signed(64'sh0) : $signed(_GEN_135); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_137 = 4'h4 == _T_9 ? $signed(regsB_1_re) : $signed(_GEN_136); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_138 = 4'h5 == _T_9 ? $signed(64'sh0) : $signed(_GEN_137); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_139 = 4'h6 == _T_9 ? $signed(64'sh0) : $signed(_GEN_138); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_140 = 4'h7 == _T_9 ? $signed(64'sh0) : $signed(_GEN_139); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_141 = 4'h8 == _T_9 ? $signed(regsB_2_re) : $signed(_GEN_140); // @[Matrix_Mul_V1.scala 162:{19,19}]
  PE PE ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_clock),
    .io_reset(PE_io_reset),
    .io_in_x_re(PE_io_in_x_re),
    .io_in_x_im(PE_io_in_x_im),
    .io_in_y_re(PE_io_in_y_re),
    .io_in_y_im(PE_io_in_y_im),
    .io_out_pe_re(PE_io_out_pe_re),
    .io_out_pe_im(PE_io_out_pe_im),
    .io_out_x_re(PE_io_out_x_re),
    .io_out_x_im(PE_io_out_x_im),
    .io_out_y_re(PE_io_out_y_re),
    .io_out_y_im(PE_io_out_y_im)
  );
  PE PE_1 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_1_clock),
    .io_reset(PE_1_io_reset),
    .io_in_x_re(PE_1_io_in_x_re),
    .io_in_x_im(PE_1_io_in_x_im),
    .io_in_y_re(PE_1_io_in_y_re),
    .io_in_y_im(PE_1_io_in_y_im),
    .io_out_pe_re(PE_1_io_out_pe_re),
    .io_out_pe_im(PE_1_io_out_pe_im),
    .io_out_x_re(PE_1_io_out_x_re),
    .io_out_x_im(PE_1_io_out_x_im),
    .io_out_y_re(PE_1_io_out_y_re),
    .io_out_y_im(PE_1_io_out_y_im)
  );
  PE PE_2 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_2_clock),
    .io_reset(PE_2_io_reset),
    .io_in_x_re(PE_2_io_in_x_re),
    .io_in_x_im(PE_2_io_in_x_im),
    .io_in_y_re(PE_2_io_in_y_re),
    .io_in_y_im(PE_2_io_in_y_im),
    .io_out_pe_re(PE_2_io_out_pe_re),
    .io_out_pe_im(PE_2_io_out_pe_im),
    .io_out_x_re(PE_2_io_out_x_re),
    .io_out_x_im(PE_2_io_out_x_im),
    .io_out_y_re(PE_2_io_out_y_re),
    .io_out_y_im(PE_2_io_out_y_im)
  );
  PE PE_3 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_3_clock),
    .io_reset(PE_3_io_reset),
    .io_in_x_re(PE_3_io_in_x_re),
    .io_in_x_im(PE_3_io_in_x_im),
    .io_in_y_re(PE_3_io_in_y_re),
    .io_in_y_im(PE_3_io_in_y_im),
    .io_out_pe_re(PE_3_io_out_pe_re),
    .io_out_pe_im(PE_3_io_out_pe_im),
    .io_out_x_re(PE_3_io_out_x_re),
    .io_out_x_im(PE_3_io_out_x_im),
    .io_out_y_re(PE_3_io_out_y_re),
    .io_out_y_im(PE_3_io_out_y_im)
  );
  PE PE_4 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_4_clock),
    .io_reset(PE_4_io_reset),
    .io_in_x_re(PE_4_io_in_x_re),
    .io_in_x_im(PE_4_io_in_x_im),
    .io_in_y_re(PE_4_io_in_y_re),
    .io_in_y_im(PE_4_io_in_y_im),
    .io_out_pe_re(PE_4_io_out_pe_re),
    .io_out_pe_im(PE_4_io_out_pe_im),
    .io_out_x_re(PE_4_io_out_x_re),
    .io_out_x_im(PE_4_io_out_x_im),
    .io_out_y_re(PE_4_io_out_y_re),
    .io_out_y_im(PE_4_io_out_y_im)
  );
  PE PE_5 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_5_clock),
    .io_reset(PE_5_io_reset),
    .io_in_x_re(PE_5_io_in_x_re),
    .io_in_x_im(PE_5_io_in_x_im),
    .io_in_y_re(PE_5_io_in_y_re),
    .io_in_y_im(PE_5_io_in_y_im),
    .io_out_pe_re(PE_5_io_out_pe_re),
    .io_out_pe_im(PE_5_io_out_pe_im),
    .io_out_x_re(PE_5_io_out_x_re),
    .io_out_x_im(PE_5_io_out_x_im),
    .io_out_y_re(PE_5_io_out_y_re),
    .io_out_y_im(PE_5_io_out_y_im)
  );
  PE PE_6 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_6_clock),
    .io_reset(PE_6_io_reset),
    .io_in_x_re(PE_6_io_in_x_re),
    .io_in_x_im(PE_6_io_in_x_im),
    .io_in_y_re(PE_6_io_in_y_re),
    .io_in_y_im(PE_6_io_in_y_im),
    .io_out_pe_re(PE_6_io_out_pe_re),
    .io_out_pe_im(PE_6_io_out_pe_im),
    .io_out_x_re(PE_6_io_out_x_re),
    .io_out_x_im(PE_6_io_out_x_im),
    .io_out_y_re(PE_6_io_out_y_re),
    .io_out_y_im(PE_6_io_out_y_im)
  );
  PE PE_7 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_7_clock),
    .io_reset(PE_7_io_reset),
    .io_in_x_re(PE_7_io_in_x_re),
    .io_in_x_im(PE_7_io_in_x_im),
    .io_in_y_re(PE_7_io_in_y_re),
    .io_in_y_im(PE_7_io_in_y_im),
    .io_out_pe_re(PE_7_io_out_pe_re),
    .io_out_pe_im(PE_7_io_out_pe_im),
    .io_out_x_re(PE_7_io_out_x_re),
    .io_out_x_im(PE_7_io_out_x_im),
    .io_out_y_re(PE_7_io_out_y_re),
    .io_out_y_im(PE_7_io_out_y_im)
  );
  PE PE_8 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_8_clock),
    .io_reset(PE_8_io_reset),
    .io_in_x_re(PE_8_io_in_x_re),
    .io_in_x_im(PE_8_io_in_x_im),
    .io_in_y_re(PE_8_io_in_y_re),
    .io_in_y_im(PE_8_io_in_y_im),
    .io_out_pe_re(PE_8_io_out_pe_re),
    .io_out_pe_im(PE_8_io_out_pe_im),
    .io_out_x_re(PE_8_io_out_x_re),
    .io_out_x_im(PE_8_io_out_x_im),
    .io_out_y_re(PE_8_io_out_y_re),
    .io_out_y_im(PE_8_io_out_y_im)
  );
  assign io_matrixC_0_re = PE_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_0_im = PE_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_1_re = PE_1_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_1_im = PE_1_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_2_re = PE_2_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_2_im = PE_2_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_3_re = PE_3_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_3_im = PE_3_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_4_re = PE_4_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_4_im = PE_4_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_5_re = PE_5_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_5_im = PE_5_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_6_re = PE_6_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_6_im = PE_6_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_7_re = PE_7_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_7_im = PE_7_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_8_re = PE_8_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_8_im = PE_8_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_valid = input_point >= 4'h5; // @[Matrix_Mul_V1.scala 188:20]
  assign PE_clock = clock;
  assign PE_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_io_in_x_re = input_point < 4'h3 ? $signed(_GEN_45) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_io_in_x_im = input_point < 4'h3 ? $signed(_GEN_36) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_io_in_y_re = _T ? $signed(_GEN_105) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_io_in_y_im = _T ? $signed(_GEN_96) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_1_clock = clock;
  assign PE_1_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_1_io_in_x_re = PE_io_out_x_re; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_1_io_in_x_im = PE_io_out_x_im; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_1_io_in_y_re = _T ? $signed(_GEN_123) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_1_io_in_y_im = _T ? $signed(_GEN_114) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_2_clock = clock;
  assign PE_2_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_2_io_in_x_re = PE_1_io_out_x_re; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_2_io_in_x_im = PE_1_io_out_x_im; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_2_io_in_y_re = _T ? $signed(_GEN_141) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_2_io_in_y_im = _T ? $signed(_GEN_132) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_3_clock = clock;
  assign PE_3_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_3_io_in_x_re = input_point < 4'h3 ? $signed(_GEN_63) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_3_io_in_x_im = input_point < 4'h3 ? $signed(_GEN_54) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_3_io_in_y_re = PE_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_3_io_in_y_im = PE_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_4_clock = clock;
  assign PE_4_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_4_io_in_x_re = PE_3_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_4_io_in_x_im = PE_3_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_4_io_in_y_re = PE_1_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_4_io_in_y_im = PE_1_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_5_clock = clock;
  assign PE_5_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_5_io_in_x_re = PE_4_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_5_io_in_x_im = PE_4_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_5_io_in_y_re = PE_2_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_5_io_in_y_im = PE_2_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_6_clock = clock;
  assign PE_6_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_6_io_in_x_re = input_point < 4'h3 ? $signed(_GEN_81) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_6_io_in_x_im = input_point < 4'h3 ? $signed(_GEN_72) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_6_io_in_y_re = PE_3_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_6_io_in_y_im = PE_3_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_7_clock = clock;
  assign PE_7_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_7_io_in_x_re = PE_6_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_7_io_in_x_im = PE_6_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_7_io_in_y_re = PE_4_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_7_io_in_y_im = PE_4_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_8_clock = clock;
  assign PE_8_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_8_io_in_x_re = PE_7_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_8_io_in_x_im = PE_7_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_8_io_in_y_re = PE_5_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_8_io_in_y_im = PE_5_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  always @(posedge clock) begin
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_0_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_0_re <= io_matrixA_0_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_0_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_0_im <= io_matrixA_0_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_1_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_1_re <= io_matrixA_1_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_1_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_1_im <= io_matrixA_1_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_2_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_2_re <= io_matrixA_2_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_2_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_2_im <= io_matrixA_2_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_0_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_0_re <= io_matrixB_0_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_0_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_0_im <= io_matrixB_0_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_1_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_1_re <= io_matrixB_1_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_1_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_1_im <= io_matrixB_1_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_2_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_2_re <= io_matrixB_2_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_2_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_2_im <= io_matrixB_2_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      input_point <= 4'h0; // @[Matrix_Mul_V1.scala 99:17]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      input_point <= 4'h0; // @[Matrix_Mul_V1.scala 108:17]
    end else begin
      input_point <= _input_point_T_1; // @[Matrix_Mul_V1.scala 116:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regsA_0_re = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regsA_0_im = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  regsA_1_re = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  regsA_1_im = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  regsA_2_re = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  regsA_2_im = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  regsB_0_re = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  regsB_0_im = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  regsB_1_re = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  regsB_1_im = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  regsB_2_re = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  regsB_2_im = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  input_point = _RAND_12[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ComplexSub(
  input  [63:0] io_op1_re,
  input  [63:0] io_op1_im,
  input  [63:0] io_op2_re,
  input  [63:0] io_op2_im,
  output [63:0] io_res_re,
  output [63:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) - $signed(io_op2_re); // @[Complex_Operater.scala 22:26]
  assign io_res_im = $signed(io_op1_im) - $signed(io_op2_im); // @[Complex_Operater.scala 23:26]
endmodule
module cholesky_comp_unit(
  input         clock,
  input         reset,
  input         io_reset,
  input         io_ready,
  input  [63:0] io_matrixIn_0_re,
  input  [63:0] io_matrixIn_0_im,
  input  [63:0] io_matrixIn_1_re,
  input  [63:0] io_matrixIn_1_im,
  input  [63:0] io_matrixIn_2_re,
  input  [63:0] io_matrixIn_2_im,
  input  [63:0] io_matrixIn_3_re,
  input  [63:0] io_matrixIn_3_im,
  input  [63:0] io_matrixIn_4_re,
  input  [63:0] io_matrixIn_4_im,
  input  [63:0] io_matrixIn_5_re,
  input  [63:0] io_matrixIn_5_im,
  input  [63:0] io_matrixIn_6_re,
  input  [63:0] io_matrixIn_6_im,
  input  [63:0] io_matrixIn_7_re,
  input  [63:0] io_matrixIn_7_im,
  input  [63:0] io_matrixIn_8_re,
  input  [63:0] io_matrixIn_8_im,
  input  [63:0] io_matrixIn_9_re,
  input  [63:0] io_matrixIn_9_im,
  input  [63:0] io_matrixIn_10_re,
  input  [63:0] io_matrixIn_10_im,
  input  [63:0] io_matrixIn_11_re,
  input  [63:0] io_matrixIn_11_im,
  input  [63:0] io_matrixIn_12_re,
  input  [63:0] io_matrixIn_12_im,
  input  [63:0] io_matrixIn_13_re,
  input  [63:0] io_matrixIn_13_im,
  input  [63:0] io_matrixIn_14_re,
  input  [63:0] io_matrixIn_14_im,
  input  [63:0] io_matrixIn_15_re,
  input  [63:0] io_matrixIn_15_im,
  output [63:0] io_matrixOut_0_re,
  output [63:0] io_matrixOut_0_im,
  output [63:0] io_matrixOut_1_re,
  output [63:0] io_matrixOut_1_im,
  output [63:0] io_matrixOut_2_re,
  output [63:0] io_matrixOut_2_im,
  output [63:0] io_matrixOut_3_re,
  output [63:0] io_matrixOut_3_im,
  output [63:0] io_matrixOut_4_re,
  output [63:0] io_matrixOut_4_im,
  output [63:0] io_matrixOut_5_re,
  output [63:0] io_matrixOut_5_im,
  output [63:0] io_matrixOut_6_re,
  output [63:0] io_matrixOut_6_im,
  output [63:0] io_matrixOut_7_re,
  output [63:0] io_matrixOut_7_im,
  output [63:0] io_matrixOut_8_re,
  output [63:0] io_matrixOut_8_im,
  output [63:0] io_matrixOut_9_re,
  output [63:0] io_matrixOut_9_im,
  output [63:0] io_matrixOut_10_re,
  output [63:0] io_matrixOut_10_im,
  output [63:0] io_matrixOut_11_re,
  output [63:0] io_matrixOut_11_im,
  output [63:0] io_matrixOut_12_re,
  output [63:0] io_matrixOut_12_im,
  output [63:0] io_matrixOut_13_re,
  output [63:0] io_matrixOut_13_im,
  output [63:0] io_matrixOut_14_re,
  output [63:0] io_matrixOut_14_im,
  output [63:0] io_matrixOut_15_re,
  output [63:0] io_matrixOut_15_im,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  wire  complex_square_root_unit_clock; // @[Cholesky_V1.scala 30:68]
  wire  complex_square_root_unit_reset; // @[Cholesky_V1.scala 30:68]
  wire [63:0] complex_square_root_unit_io_op_re; // @[Cholesky_V1.scala 30:68]
  wire [63:0] complex_square_root_unit_io_op_im; // @[Cholesky_V1.scala 30:68]
  wire [63:0] complex_square_root_unit_io_res_re; // @[Cholesky_V1.scala 30:68]
  wire [63:0] complex_square_root_unit_io_res_im; // @[Cholesky_V1.scala 30:68]
  wire  complex_divide_unit_clock; // @[Cholesky_V1.scala 31:58]
  wire  complex_divide_unit_reset; // @[Cholesky_V1.scala 31:58]
  wire [63:0] complex_divide_unit_io_op2_re; // @[Cholesky_V1.scala 31:58]
  wire [63:0] complex_divide_unit_io_op2_im; // @[Cholesky_V1.scala 31:58]
  wire [63:0] complex_divide_unit_io_res_re; // @[Cholesky_V1.scala 31:58]
  wire [63:0] complex_divide_unit_io_res_im; // @[Cholesky_V1.scala 31:58]
  wire  matirx_mul_unit_clock; // @[Cholesky_V1.scala 32:46]
  wire  matirx_mul_unit_io_reset; // @[Cholesky_V1.scala 32:46]
  wire  matirx_mul_unit_io_ready; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixA_0_re; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixA_0_im; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixA_1_re; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixA_1_im; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixA_2_re; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixA_2_im; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixB_0_re; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixB_0_im; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixB_1_re; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixB_1_im; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixB_2_re; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixB_2_im; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_0_re; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_0_im; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_1_re; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_1_im; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_2_re; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_2_im; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_3_re; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_3_im; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_4_re; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_4_im; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_5_re; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_5_im; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_6_re; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_6_im; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_7_re; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_7_im; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_8_re; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matirx_mul_unit_io_matrixC_8_im; // @[Cholesky_V1.scala 32:46]
  wire  matirx_mul_unit_io_valid; // @[Cholesky_V1.scala 32:46]
  wire [63:0] matrix_comp_reg_4_mul_io_op1_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] matrix_comp_reg_4_mul_io_op1_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] matrix_comp_reg_4_mul_io_op2_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] matrix_comp_reg_4_mul_io_op2_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] matrix_comp_reg_4_mul_io_res_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] matrix_comp_reg_4_mul_io_res_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] matrix_comp_reg_8_mul_io_op1_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] matrix_comp_reg_8_mul_io_op1_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] matrix_comp_reg_8_mul_io_op2_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] matrix_comp_reg_8_mul_io_op2_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] matrix_comp_reg_8_mul_io_res_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] matrix_comp_reg_8_mul_io_res_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] matrix_comp_reg_12_mul_io_op1_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] matrix_comp_reg_12_mul_io_op1_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] matrix_comp_reg_12_mul_io_op2_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] matrix_comp_reg_12_mul_io_op2_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] matrix_comp_reg_12_mul_io_res_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] matrix_comp_reg_12_mul_io_res_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_5_sub_io_op1_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_5_sub_io_op1_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_5_sub_io_op2_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_5_sub_io_op2_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_5_sub_io_res_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_5_sub_io_res_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_6_sub_io_op1_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_6_sub_io_op1_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_6_sub_io_op2_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_6_sub_io_op2_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_6_sub_io_res_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_6_sub_io_res_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_7_sub_io_op1_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_7_sub_io_op1_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_7_sub_io_op2_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_7_sub_io_op2_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_7_sub_io_res_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_7_sub_io_res_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_9_sub_io_op1_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_9_sub_io_op1_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_9_sub_io_op2_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_9_sub_io_op2_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_9_sub_io_res_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_9_sub_io_res_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_10_sub_io_op1_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_10_sub_io_op1_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_10_sub_io_op2_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_10_sub_io_op2_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_10_sub_io_res_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_10_sub_io_res_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_11_sub_io_op1_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_11_sub_io_op1_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_11_sub_io_op2_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_11_sub_io_op2_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_11_sub_io_res_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_11_sub_io_res_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_13_sub_io_op1_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_13_sub_io_op1_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_13_sub_io_op2_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_13_sub_io_op2_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_13_sub_io_res_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_13_sub_io_res_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_14_sub_io_op1_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_14_sub_io_op1_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_14_sub_io_op2_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_14_sub_io_op2_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_14_sub_io_res_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_14_sub_io_res_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_15_sub_io_op1_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_15_sub_io_op1_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_15_sub_io_op2_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_15_sub_io_op2_im; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_15_sub_io_res_re; // @[Complex_Operater.scala 29:21]
  wire [63:0] io_matrixOut_15_sub_io_res_im; // @[Complex_Operater.scala 29:21]
  reg [63:0] matrix_comp_reg_0_re; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_0_im; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_1_re; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_1_im; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_2_re; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_2_im; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_3_re; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_3_im; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_4_re; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_4_im; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_5_re; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_5_im; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_6_re; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_6_im; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_7_re; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_7_im; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_8_re; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_8_im; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_9_re; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_9_im; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_10_re; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_10_im; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_11_re; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_11_im; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_12_re; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_12_im; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_13_re; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_13_im; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_14_re; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_14_im; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_15_re; // @[Cholesky_V1.scala 23:42]
  reg [63:0] matrix_comp_reg_15_im; // @[Cholesky_V1.scala 23:42]
  reg [7:0] status; // @[Cholesky_V1.scala 24:29]
  wire [7:0] _status_T_1 = status + 8'h1; // @[Cholesky_V1.scala 59:24]
  wire [7:0] _GEN_0 = matirx_mul_unit_io_valid ? _status_T_1 : status; // @[Cholesky_V1.scala 81:38 82:16 24:29]
  wire [7:0] _GEN_2 = status == 8'h50 ? _GEN_0 : status; // @[Cholesky_V1.scala 24:29 79:55]
  wire [7:0] _GEN_10 = status == 8'h4f ? _status_T_1 : _GEN_2; // @[Cholesky_V1.scala 74:55 78:14]
  wire [63:0] _GEN_11 = status == 8'h4e ? $signed(matrix_comp_reg_4_mul_io_res_im) : $signed(matrix_comp_reg_4_im); // @[Cholesky_V1.scala 23:42 68:55 71:42]
  wire [63:0] _GEN_12 = status == 8'h4e ? $signed(matrix_comp_reg_4_mul_io_res_re) : $signed(matrix_comp_reg_4_re); // @[Cholesky_V1.scala 23:42 68:55 71:42]
  wire [63:0] _GEN_13 = status == 8'h4e ? $signed(matrix_comp_reg_8_mul_io_res_im) : $signed(matrix_comp_reg_8_im); // @[Cholesky_V1.scala 23:42 68:55 71:42]
  wire [63:0] _GEN_14 = status == 8'h4e ? $signed(matrix_comp_reg_8_mul_io_res_re) : $signed(matrix_comp_reg_8_re); // @[Cholesky_V1.scala 23:42 68:55 71:42]
  wire [63:0] _GEN_15 = status == 8'h4e ? $signed(matrix_comp_reg_12_mul_io_res_im) : $signed(matrix_comp_reg_12_im); // @[Cholesky_V1.scala 23:42 68:55 71:42]
  wire [63:0] _GEN_16 = status == 8'h4e ? $signed(matrix_comp_reg_12_mul_io_res_re) : $signed(matrix_comp_reg_12_re); // @[Cholesky_V1.scala 23:42 68:55 71:42]
  wire [7:0] _GEN_17 = status == 8'h4e ? _status_T_1 : _GEN_10; // @[Cholesky_V1.scala 68:55 73:14]
  wire [63:0] _GEN_25 = status <= 8'h4d ? $signed(matrix_comp_reg_0_im) : $signed(64'sh100000000); // @[Cholesky_V1.scala 37:33 64:54 66:34]
  wire [63:0] _GEN_26 = status <= 8'h4d ? $signed(matrix_comp_reg_0_re) : $signed(64'sh100000000); // @[Cholesky_V1.scala 36:33 64:54 66:34]
  wire [7:0] _GEN_27 = status <= 8'h4d ? _status_T_1 : _GEN_17; // @[Cholesky_V1.scala 64:54 67:14]
  wire [63:0] _GEN_28 = status <= 8'h4d ? $signed(matrix_comp_reg_4_im) : $signed(_GEN_11); // @[Cholesky_V1.scala 23:42 64:54]
  wire [63:0] _GEN_29 = status <= 8'h4d ? $signed(matrix_comp_reg_4_re) : $signed(_GEN_12); // @[Cholesky_V1.scala 23:42 64:54]
  wire [63:0] _GEN_30 = status <= 8'h4d ? $signed(matrix_comp_reg_8_im) : $signed(_GEN_13); // @[Cholesky_V1.scala 23:42 64:54]
  wire [63:0] _GEN_31 = status <= 8'h4d ? $signed(matrix_comp_reg_8_re) : $signed(_GEN_14); // @[Cholesky_V1.scala 23:42 64:54]
  wire [63:0] _GEN_32 = status <= 8'h4d ? $signed(matrix_comp_reg_12_im) : $signed(_GEN_15); // @[Cholesky_V1.scala 23:42 64:54]
  wire [63:0] _GEN_33 = status <= 8'h4d ? $signed(matrix_comp_reg_12_re) : $signed(_GEN_16); // @[Cholesky_V1.scala 23:42 64:54]
  wire [7:0] _GEN_43 = status == 8'h20 ? _status_T_1 : _GEN_27; // @[Cholesky_V1.scala 60:55 63:14]
  wire [63:0] _GEN_44 = status == 8'h20 ? $signed(64'sh100000000) : $signed(_GEN_25); // @[Cholesky_V1.scala 37:33 60:55]
  wire [63:0] _GEN_45 = status == 8'h20 ? $signed(64'sh100000000) : $signed(_GEN_26); // @[Cholesky_V1.scala 36:33 60:55]
  wire [63:0] _GEN_64 = status <= 8'h1f ? $signed(64'sh100000000) : $signed(_GEN_44); // @[Cholesky_V1.scala 37:33 56:48]
  wire [63:0] _GEN_65 = status <= 8'h1f ? $signed(64'sh100000000) : $signed(_GEN_45); // @[Cholesky_V1.scala 36:33 56:48]
  wire [63:0] _GEN_114 = io_ready ? $signed(64'sh100000000) : $signed(_GEN_64); // @[Cholesky_V1.scala 50:24 37:33]
  wire [63:0] _GEN_115 = io_ready ? $signed(64'sh100000000) : $signed(_GEN_65); // @[Cholesky_V1.scala 50:24 36:33]
  cordic_complex_square_root complex_square_root_unit ( // @[Cholesky_V1.scala 30:68]
    .clock(complex_square_root_unit_clock),
    .reset(complex_square_root_unit_reset),
    .io_op_re(complex_square_root_unit_io_op_re),
    .io_op_im(complex_square_root_unit_io_op_im),
    .io_res_re(complex_square_root_unit_io_res_re),
    .io_res_im(complex_square_root_unit_io_res_im)
  );
  cordic_complex_divide complex_divide_unit ( // @[Cholesky_V1.scala 31:58]
    .clock(complex_divide_unit_clock),
    .reset(complex_divide_unit_reset),
    .io_op2_re(complex_divide_unit_io_op2_re),
    .io_op2_im(complex_divide_unit_io_op2_im),
    .io_res_re(complex_divide_unit_io_res_re),
    .io_res_im(complex_divide_unit_io_res_im)
  );
  matrix_mul_v1_1 matirx_mul_unit ( // @[Cholesky_V1.scala 32:46]
    .clock(matirx_mul_unit_clock),
    .io_reset(matirx_mul_unit_io_reset),
    .io_ready(matirx_mul_unit_io_ready),
    .io_matrixA_0_re(matirx_mul_unit_io_matrixA_0_re),
    .io_matrixA_0_im(matirx_mul_unit_io_matrixA_0_im),
    .io_matrixA_1_re(matirx_mul_unit_io_matrixA_1_re),
    .io_matrixA_1_im(matirx_mul_unit_io_matrixA_1_im),
    .io_matrixA_2_re(matirx_mul_unit_io_matrixA_2_re),
    .io_matrixA_2_im(matirx_mul_unit_io_matrixA_2_im),
    .io_matrixB_0_re(matirx_mul_unit_io_matrixB_0_re),
    .io_matrixB_0_im(matirx_mul_unit_io_matrixB_0_im),
    .io_matrixB_1_re(matirx_mul_unit_io_matrixB_1_re),
    .io_matrixB_1_im(matirx_mul_unit_io_matrixB_1_im),
    .io_matrixB_2_re(matirx_mul_unit_io_matrixB_2_re),
    .io_matrixB_2_im(matirx_mul_unit_io_matrixB_2_im),
    .io_matrixC_0_re(matirx_mul_unit_io_matrixC_0_re),
    .io_matrixC_0_im(matirx_mul_unit_io_matrixC_0_im),
    .io_matrixC_1_re(matirx_mul_unit_io_matrixC_1_re),
    .io_matrixC_1_im(matirx_mul_unit_io_matrixC_1_im),
    .io_matrixC_2_re(matirx_mul_unit_io_matrixC_2_re),
    .io_matrixC_2_im(matirx_mul_unit_io_matrixC_2_im),
    .io_matrixC_3_re(matirx_mul_unit_io_matrixC_3_re),
    .io_matrixC_3_im(matirx_mul_unit_io_matrixC_3_im),
    .io_matrixC_4_re(matirx_mul_unit_io_matrixC_4_re),
    .io_matrixC_4_im(matirx_mul_unit_io_matrixC_4_im),
    .io_matrixC_5_re(matirx_mul_unit_io_matrixC_5_re),
    .io_matrixC_5_im(matirx_mul_unit_io_matrixC_5_im),
    .io_matrixC_6_re(matirx_mul_unit_io_matrixC_6_re),
    .io_matrixC_6_im(matirx_mul_unit_io_matrixC_6_im),
    .io_matrixC_7_re(matirx_mul_unit_io_matrixC_7_re),
    .io_matrixC_7_im(matirx_mul_unit_io_matrixC_7_im),
    .io_matrixC_8_re(matirx_mul_unit_io_matrixC_8_re),
    .io_matrixC_8_im(matirx_mul_unit_io_matrixC_8_im),
    .io_valid(matirx_mul_unit_io_valid)
  );
  ComplexMul matrix_comp_reg_4_mul ( // @[Complex_Operater.scala 47:21]
    .io_op1_re(matrix_comp_reg_4_mul_io_op1_re),
    .io_op1_im(matrix_comp_reg_4_mul_io_op1_im),
    .io_op2_re(matrix_comp_reg_4_mul_io_op2_re),
    .io_op2_im(matrix_comp_reg_4_mul_io_op2_im),
    .io_res_re(matrix_comp_reg_4_mul_io_res_re),
    .io_res_im(matrix_comp_reg_4_mul_io_res_im)
  );
  ComplexMul matrix_comp_reg_8_mul ( // @[Complex_Operater.scala 47:21]
    .io_op1_re(matrix_comp_reg_8_mul_io_op1_re),
    .io_op1_im(matrix_comp_reg_8_mul_io_op1_im),
    .io_op2_re(matrix_comp_reg_8_mul_io_op2_re),
    .io_op2_im(matrix_comp_reg_8_mul_io_op2_im),
    .io_res_re(matrix_comp_reg_8_mul_io_res_re),
    .io_res_im(matrix_comp_reg_8_mul_io_res_im)
  );
  ComplexMul matrix_comp_reg_12_mul ( // @[Complex_Operater.scala 47:21]
    .io_op1_re(matrix_comp_reg_12_mul_io_op1_re),
    .io_op1_im(matrix_comp_reg_12_mul_io_op1_im),
    .io_op2_re(matrix_comp_reg_12_mul_io_op2_re),
    .io_op2_im(matrix_comp_reg_12_mul_io_op2_im),
    .io_res_re(matrix_comp_reg_12_mul_io_res_re),
    .io_res_im(matrix_comp_reg_12_mul_io_res_im)
  );
  ComplexSub io_matrixOut_5_sub ( // @[Complex_Operater.scala 29:21]
    .io_op1_re(io_matrixOut_5_sub_io_op1_re),
    .io_op1_im(io_matrixOut_5_sub_io_op1_im),
    .io_op2_re(io_matrixOut_5_sub_io_op2_re),
    .io_op2_im(io_matrixOut_5_sub_io_op2_im),
    .io_res_re(io_matrixOut_5_sub_io_res_re),
    .io_res_im(io_matrixOut_5_sub_io_res_im)
  );
  ComplexSub io_matrixOut_6_sub ( // @[Complex_Operater.scala 29:21]
    .io_op1_re(io_matrixOut_6_sub_io_op1_re),
    .io_op1_im(io_matrixOut_6_sub_io_op1_im),
    .io_op2_re(io_matrixOut_6_sub_io_op2_re),
    .io_op2_im(io_matrixOut_6_sub_io_op2_im),
    .io_res_re(io_matrixOut_6_sub_io_res_re),
    .io_res_im(io_matrixOut_6_sub_io_res_im)
  );
  ComplexSub io_matrixOut_7_sub ( // @[Complex_Operater.scala 29:21]
    .io_op1_re(io_matrixOut_7_sub_io_op1_re),
    .io_op1_im(io_matrixOut_7_sub_io_op1_im),
    .io_op2_re(io_matrixOut_7_sub_io_op2_re),
    .io_op2_im(io_matrixOut_7_sub_io_op2_im),
    .io_res_re(io_matrixOut_7_sub_io_res_re),
    .io_res_im(io_matrixOut_7_sub_io_res_im)
  );
  ComplexSub io_matrixOut_9_sub ( // @[Complex_Operater.scala 29:21]
    .io_op1_re(io_matrixOut_9_sub_io_op1_re),
    .io_op1_im(io_matrixOut_9_sub_io_op1_im),
    .io_op2_re(io_matrixOut_9_sub_io_op2_re),
    .io_op2_im(io_matrixOut_9_sub_io_op2_im),
    .io_res_re(io_matrixOut_9_sub_io_res_re),
    .io_res_im(io_matrixOut_9_sub_io_res_im)
  );
  ComplexSub io_matrixOut_10_sub ( // @[Complex_Operater.scala 29:21]
    .io_op1_re(io_matrixOut_10_sub_io_op1_re),
    .io_op1_im(io_matrixOut_10_sub_io_op1_im),
    .io_op2_re(io_matrixOut_10_sub_io_op2_re),
    .io_op2_im(io_matrixOut_10_sub_io_op2_im),
    .io_res_re(io_matrixOut_10_sub_io_res_re),
    .io_res_im(io_matrixOut_10_sub_io_res_im)
  );
  ComplexSub io_matrixOut_11_sub ( // @[Complex_Operater.scala 29:21]
    .io_op1_re(io_matrixOut_11_sub_io_op1_re),
    .io_op1_im(io_matrixOut_11_sub_io_op1_im),
    .io_op2_re(io_matrixOut_11_sub_io_op2_re),
    .io_op2_im(io_matrixOut_11_sub_io_op2_im),
    .io_res_re(io_matrixOut_11_sub_io_res_re),
    .io_res_im(io_matrixOut_11_sub_io_res_im)
  );
  ComplexSub io_matrixOut_13_sub ( // @[Complex_Operater.scala 29:21]
    .io_op1_re(io_matrixOut_13_sub_io_op1_re),
    .io_op1_im(io_matrixOut_13_sub_io_op1_im),
    .io_op2_re(io_matrixOut_13_sub_io_op2_re),
    .io_op2_im(io_matrixOut_13_sub_io_op2_im),
    .io_res_re(io_matrixOut_13_sub_io_res_re),
    .io_res_im(io_matrixOut_13_sub_io_res_im)
  );
  ComplexSub io_matrixOut_14_sub ( // @[Complex_Operater.scala 29:21]
    .io_op1_re(io_matrixOut_14_sub_io_op1_re),
    .io_op1_im(io_matrixOut_14_sub_io_op1_im),
    .io_op2_re(io_matrixOut_14_sub_io_op2_re),
    .io_op2_im(io_matrixOut_14_sub_io_op2_im),
    .io_res_re(io_matrixOut_14_sub_io_res_re),
    .io_res_im(io_matrixOut_14_sub_io_res_im)
  );
  ComplexSub io_matrixOut_15_sub ( // @[Complex_Operater.scala 29:21]
    .io_op1_re(io_matrixOut_15_sub_io_op1_re),
    .io_op1_im(io_matrixOut_15_sub_io_op1_im),
    .io_op2_re(io_matrixOut_15_sub_io_op2_re),
    .io_op2_im(io_matrixOut_15_sub_io_op2_im),
    .io_res_re(io_matrixOut_15_sub_io_res_re),
    .io_res_im(io_matrixOut_15_sub_io_res_im)
  );
  assign io_matrixOut_0_re = matrix_comp_reg_0_re; // @[Cholesky_V1.scala 93:16]
  assign io_matrixOut_0_im = matrix_comp_reg_0_im; // @[Cholesky_V1.scala 93:16]
  assign io_matrixOut_1_re = matrix_comp_reg_1_re; // @[Cholesky_V1.scala 93:16]
  assign io_matrixOut_1_im = matrix_comp_reg_1_im; // @[Cholesky_V1.scala 93:16]
  assign io_matrixOut_2_re = matrix_comp_reg_2_re; // @[Cholesky_V1.scala 93:16]
  assign io_matrixOut_2_im = matrix_comp_reg_2_im; // @[Cholesky_V1.scala 93:16]
  assign io_matrixOut_3_re = matrix_comp_reg_3_re; // @[Cholesky_V1.scala 93:16]
  assign io_matrixOut_3_im = matrix_comp_reg_3_im; // @[Cholesky_V1.scala 93:16]
  assign io_matrixOut_4_re = matrix_comp_reg_4_re; // @[Cholesky_V1.scala 93:16]
  assign io_matrixOut_4_im = matrix_comp_reg_4_im; // @[Cholesky_V1.scala 93:16]
  assign io_matrixOut_5_re = io_matrixOut_5_sub_io_res_re; // @[Cholesky_V1.scala 96:43]
  assign io_matrixOut_5_im = io_matrixOut_5_sub_io_res_im; // @[Cholesky_V1.scala 96:43]
  assign io_matrixOut_6_re = io_matrixOut_6_sub_io_res_re; // @[Cholesky_V1.scala 96:43]
  assign io_matrixOut_6_im = io_matrixOut_6_sub_io_res_im; // @[Cholesky_V1.scala 96:43]
  assign io_matrixOut_7_re = io_matrixOut_7_sub_io_res_re; // @[Cholesky_V1.scala 96:43]
  assign io_matrixOut_7_im = io_matrixOut_7_sub_io_res_im; // @[Cholesky_V1.scala 96:43]
  assign io_matrixOut_8_re = matrix_comp_reg_8_re; // @[Cholesky_V1.scala 93:16]
  assign io_matrixOut_8_im = matrix_comp_reg_8_im; // @[Cholesky_V1.scala 93:16]
  assign io_matrixOut_9_re = io_matrixOut_9_sub_io_res_re; // @[Cholesky_V1.scala 96:43]
  assign io_matrixOut_9_im = io_matrixOut_9_sub_io_res_im; // @[Cholesky_V1.scala 96:43]
  assign io_matrixOut_10_re = io_matrixOut_10_sub_io_res_re; // @[Cholesky_V1.scala 96:43]
  assign io_matrixOut_10_im = io_matrixOut_10_sub_io_res_im; // @[Cholesky_V1.scala 96:43]
  assign io_matrixOut_11_re = io_matrixOut_11_sub_io_res_re; // @[Cholesky_V1.scala 96:43]
  assign io_matrixOut_11_im = io_matrixOut_11_sub_io_res_im; // @[Cholesky_V1.scala 96:43]
  assign io_matrixOut_12_re = matrix_comp_reg_12_re; // @[Cholesky_V1.scala 93:16]
  assign io_matrixOut_12_im = matrix_comp_reg_12_im; // @[Cholesky_V1.scala 93:16]
  assign io_matrixOut_13_re = io_matrixOut_13_sub_io_res_re; // @[Cholesky_V1.scala 96:43]
  assign io_matrixOut_13_im = io_matrixOut_13_sub_io_res_im; // @[Cholesky_V1.scala 96:43]
  assign io_matrixOut_14_re = io_matrixOut_14_sub_io_res_re; // @[Cholesky_V1.scala 96:43]
  assign io_matrixOut_14_im = io_matrixOut_14_sub_io_res_im; // @[Cholesky_V1.scala 96:43]
  assign io_matrixOut_15_re = io_matrixOut_15_sub_io_res_re; // @[Cholesky_V1.scala 96:43]
  assign io_matrixOut_15_im = io_matrixOut_15_sub_io_res_im; // @[Cholesky_V1.scala 96:43]
  assign io_valid = status > 8'h50; // @[Cholesky_V1.scala 88:15]
  assign complex_square_root_unit_clock = clock;
  assign complex_square_root_unit_reset = reset;
  assign complex_square_root_unit_io_op_re = matrix_comp_reg_0_re; // @[Cholesky_V1.scala 56:48 58:38]
  assign complex_square_root_unit_io_op_im = matrix_comp_reg_0_im; // @[Cholesky_V1.scala 56:48 58:38]
  assign complex_divide_unit_clock = clock;
  assign complex_divide_unit_reset = reset;
  assign complex_divide_unit_io_op2_re = io_reset ? $signed(64'sh100000000) : $signed(_GEN_115); // @[Cholesky_V1.scala 43:18 36:33]
  assign complex_divide_unit_io_op2_im = io_reset ? $signed(64'sh100000000) : $signed(_GEN_114); // @[Cholesky_V1.scala 43:18 37:33]
  assign matirx_mul_unit_clock = clock;
  assign matirx_mul_unit_io_reset = io_reset; // @[Cholesky_V1.scala 38:28]
  assign matirx_mul_unit_io_ready = status == 8'h4f; // @[Cholesky_V1.scala 74:23]
  assign matirx_mul_unit_io_matrixA_0_re = matrix_comp_reg_4_re; // @[Cholesky_V1.scala 25:30 27:11]
  assign matirx_mul_unit_io_matrixA_0_im = matrix_comp_reg_4_im; // @[Cholesky_V1.scala 25:30 27:11]
  assign matirx_mul_unit_io_matrixA_1_re = matrix_comp_reg_8_re; // @[Cholesky_V1.scala 25:30 27:11]
  assign matirx_mul_unit_io_matrixA_1_im = matrix_comp_reg_8_im; // @[Cholesky_V1.scala 25:30 27:11]
  assign matirx_mul_unit_io_matrixA_2_re = matrix_comp_reg_12_re; // @[Cholesky_V1.scala 25:30 27:11]
  assign matirx_mul_unit_io_matrixA_2_im = matrix_comp_reg_12_im; // @[Cholesky_V1.scala 25:30 27:11]
  assign matirx_mul_unit_io_matrixB_0_re = matrix_comp_reg_4_re; // @[Cholesky_V1.scala 25:30 27:11]
  assign matirx_mul_unit_io_matrixB_0_im = matrix_comp_reg_4_im; // @[Cholesky_V1.scala 25:30 27:11]
  assign matirx_mul_unit_io_matrixB_1_re = matrix_comp_reg_8_re; // @[Cholesky_V1.scala 25:30 27:11]
  assign matirx_mul_unit_io_matrixB_1_im = matrix_comp_reg_8_im; // @[Cholesky_V1.scala 25:30 27:11]
  assign matirx_mul_unit_io_matrixB_2_re = matrix_comp_reg_12_re; // @[Cholesky_V1.scala 25:30 27:11]
  assign matirx_mul_unit_io_matrixB_2_im = matrix_comp_reg_12_im; // @[Cholesky_V1.scala 25:30 27:11]
  assign matrix_comp_reg_4_mul_io_op1_re = matrix_comp_reg_4_re; // @[Complex_Operater.scala 48:16]
  assign matrix_comp_reg_4_mul_io_op1_im = matrix_comp_reg_4_im; // @[Complex_Operater.scala 48:16]
  assign matrix_comp_reg_4_mul_io_op2_re = complex_divide_unit_io_res_re; // @[Complex_Operater.scala 49:16]
  assign matrix_comp_reg_4_mul_io_op2_im = complex_divide_unit_io_res_im; // @[Complex_Operater.scala 49:16]
  assign matrix_comp_reg_8_mul_io_op1_re = matrix_comp_reg_8_re; // @[Complex_Operater.scala 48:16]
  assign matrix_comp_reg_8_mul_io_op1_im = matrix_comp_reg_8_im; // @[Complex_Operater.scala 48:16]
  assign matrix_comp_reg_8_mul_io_op2_re = complex_divide_unit_io_res_re; // @[Complex_Operater.scala 49:16]
  assign matrix_comp_reg_8_mul_io_op2_im = complex_divide_unit_io_res_im; // @[Complex_Operater.scala 49:16]
  assign matrix_comp_reg_12_mul_io_op1_re = matrix_comp_reg_12_re; // @[Complex_Operater.scala 48:16]
  assign matrix_comp_reg_12_mul_io_op1_im = matrix_comp_reg_12_im; // @[Complex_Operater.scala 48:16]
  assign matrix_comp_reg_12_mul_io_op2_re = complex_divide_unit_io_res_re; // @[Complex_Operater.scala 49:16]
  assign matrix_comp_reg_12_mul_io_op2_im = complex_divide_unit_io_res_im; // @[Complex_Operater.scala 49:16]
  assign io_matrixOut_5_sub_io_op1_re = matrix_comp_reg_5_re; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_5_sub_io_op1_im = matrix_comp_reg_5_im; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_5_sub_io_op2_re = matirx_mul_unit_io_matrixC_0_re; // @[Complex_Operater.scala 31:16]
  assign io_matrixOut_5_sub_io_op2_im = matirx_mul_unit_io_matrixC_0_im; // @[Complex_Operater.scala 31:16]
  assign io_matrixOut_6_sub_io_op1_re = matrix_comp_reg_6_re; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_6_sub_io_op1_im = matrix_comp_reg_6_im; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_6_sub_io_op2_re = matirx_mul_unit_io_matrixC_1_re; // @[Complex_Operater.scala 31:16]
  assign io_matrixOut_6_sub_io_op2_im = matirx_mul_unit_io_matrixC_1_im; // @[Complex_Operater.scala 31:16]
  assign io_matrixOut_7_sub_io_op1_re = matrix_comp_reg_7_re; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_7_sub_io_op1_im = matrix_comp_reg_7_im; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_7_sub_io_op2_re = matirx_mul_unit_io_matrixC_2_re; // @[Complex_Operater.scala 31:16]
  assign io_matrixOut_7_sub_io_op2_im = matirx_mul_unit_io_matrixC_2_im; // @[Complex_Operater.scala 31:16]
  assign io_matrixOut_9_sub_io_op1_re = matrix_comp_reg_9_re; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_9_sub_io_op1_im = matrix_comp_reg_9_im; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_9_sub_io_op2_re = matirx_mul_unit_io_matrixC_3_re; // @[Complex_Operater.scala 31:16]
  assign io_matrixOut_9_sub_io_op2_im = matirx_mul_unit_io_matrixC_3_im; // @[Complex_Operater.scala 31:16]
  assign io_matrixOut_10_sub_io_op1_re = matrix_comp_reg_10_re; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_10_sub_io_op1_im = matrix_comp_reg_10_im; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_10_sub_io_op2_re = matirx_mul_unit_io_matrixC_4_re; // @[Complex_Operater.scala 31:16]
  assign io_matrixOut_10_sub_io_op2_im = matirx_mul_unit_io_matrixC_4_im; // @[Complex_Operater.scala 31:16]
  assign io_matrixOut_11_sub_io_op1_re = matrix_comp_reg_11_re; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_11_sub_io_op1_im = matrix_comp_reg_11_im; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_11_sub_io_op2_re = matirx_mul_unit_io_matrixC_5_re; // @[Complex_Operater.scala 31:16]
  assign io_matrixOut_11_sub_io_op2_im = matirx_mul_unit_io_matrixC_5_im; // @[Complex_Operater.scala 31:16]
  assign io_matrixOut_13_sub_io_op1_re = matrix_comp_reg_13_re; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_13_sub_io_op1_im = matrix_comp_reg_13_im; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_13_sub_io_op2_re = matirx_mul_unit_io_matrixC_6_re; // @[Complex_Operater.scala 31:16]
  assign io_matrixOut_13_sub_io_op2_im = matirx_mul_unit_io_matrixC_6_im; // @[Complex_Operater.scala 31:16]
  assign io_matrixOut_14_sub_io_op1_re = matrix_comp_reg_14_re; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_14_sub_io_op1_im = matrix_comp_reg_14_im; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_14_sub_io_op2_re = matirx_mul_unit_io_matrixC_7_re; // @[Complex_Operater.scala 31:16]
  assign io_matrixOut_14_sub_io_op2_im = matirx_mul_unit_io_matrixC_7_im; // @[Complex_Operater.scala 31:16]
  assign io_matrixOut_15_sub_io_op1_re = matrix_comp_reg_15_re; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_15_sub_io_op1_im = matrix_comp_reg_15_im; // @[Complex_Operater.scala 30:16]
  assign io_matrixOut_15_sub_io_op2_re = matirx_mul_unit_io_matrixC_8_re; // @[Complex_Operater.scala 31:16]
  assign io_matrixOut_15_sub_io_op2_im = matirx_mul_unit_io_matrixC_8_im; // @[Complex_Operater.scala 31:16]
  always @(posedge clock) begin
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_0_re <= 64'sh0; // @[Cholesky_V1.scala 46:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_0_re <= io_matrixIn_0_re; // @[Cholesky_V1.scala 52:21]
    end else if (!(status <= 8'h1f)) begin // @[Cholesky_V1.scala 56:48]
      if (status == 8'h20) begin // @[Cholesky_V1.scala 60:55]
        matrix_comp_reg_0_re <= complex_square_root_unit_io_res_re; // @[Cholesky_V1.scala 62:26]
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_0_im <= 64'sh0; // @[Cholesky_V1.scala 47:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_0_im <= io_matrixIn_0_im; // @[Cholesky_V1.scala 52:21]
    end else if (!(status <= 8'h1f)) begin // @[Cholesky_V1.scala 56:48]
      if (status == 8'h20) begin // @[Cholesky_V1.scala 60:55]
        matrix_comp_reg_0_im <= complex_square_root_unit_io_res_im; // @[Cholesky_V1.scala 62:26]
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_1_re <= 64'sh0; // @[Cholesky_V1.scala 46:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_1_re <= io_matrixIn_1_re; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_1_im <= 64'sh0; // @[Cholesky_V1.scala 47:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_1_im <= io_matrixIn_1_im; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_2_re <= 64'sh0; // @[Cholesky_V1.scala 46:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_2_re <= io_matrixIn_2_re; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_2_im <= 64'sh0; // @[Cholesky_V1.scala 47:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_2_im <= io_matrixIn_2_im; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_3_re <= 64'sh0; // @[Cholesky_V1.scala 46:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_3_re <= io_matrixIn_3_re; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_3_im <= 64'sh0; // @[Cholesky_V1.scala 47:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_3_im <= io_matrixIn_3_im; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_4_re <= 64'sh0; // @[Cholesky_V1.scala 46:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_4_re <= io_matrixIn_4_re; // @[Cholesky_V1.scala 52:21]
    end else if (!(status <= 8'h1f)) begin // @[Cholesky_V1.scala 56:48]
      if (!(status == 8'h20)) begin // @[Cholesky_V1.scala 60:55]
        matrix_comp_reg_4_re <= _GEN_29;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_4_im <= 64'sh0; // @[Cholesky_V1.scala 47:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_4_im <= io_matrixIn_4_im; // @[Cholesky_V1.scala 52:21]
    end else if (!(status <= 8'h1f)) begin // @[Cholesky_V1.scala 56:48]
      if (!(status == 8'h20)) begin // @[Cholesky_V1.scala 60:55]
        matrix_comp_reg_4_im <= _GEN_28;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_5_re <= 64'sh0; // @[Cholesky_V1.scala 46:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_5_re <= io_matrixIn_5_re; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_5_im <= 64'sh0; // @[Cholesky_V1.scala 47:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_5_im <= io_matrixIn_5_im; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_6_re <= 64'sh0; // @[Cholesky_V1.scala 46:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_6_re <= io_matrixIn_6_re; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_6_im <= 64'sh0; // @[Cholesky_V1.scala 47:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_6_im <= io_matrixIn_6_im; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_7_re <= 64'sh0; // @[Cholesky_V1.scala 46:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_7_re <= io_matrixIn_7_re; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_7_im <= 64'sh0; // @[Cholesky_V1.scala 47:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_7_im <= io_matrixIn_7_im; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_8_re <= 64'sh0; // @[Cholesky_V1.scala 46:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_8_re <= io_matrixIn_8_re; // @[Cholesky_V1.scala 52:21]
    end else if (!(status <= 8'h1f)) begin // @[Cholesky_V1.scala 56:48]
      if (!(status == 8'h20)) begin // @[Cholesky_V1.scala 60:55]
        matrix_comp_reg_8_re <= _GEN_31;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_8_im <= 64'sh0; // @[Cholesky_V1.scala 47:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_8_im <= io_matrixIn_8_im; // @[Cholesky_V1.scala 52:21]
    end else if (!(status <= 8'h1f)) begin // @[Cholesky_V1.scala 56:48]
      if (!(status == 8'h20)) begin // @[Cholesky_V1.scala 60:55]
        matrix_comp_reg_8_im <= _GEN_30;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_9_re <= 64'sh0; // @[Cholesky_V1.scala 46:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_9_re <= io_matrixIn_9_re; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_9_im <= 64'sh0; // @[Cholesky_V1.scala 47:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_9_im <= io_matrixIn_9_im; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_10_re <= 64'sh0; // @[Cholesky_V1.scala 46:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_10_re <= io_matrixIn_10_re; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_10_im <= 64'sh0; // @[Cholesky_V1.scala 47:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_10_im <= io_matrixIn_10_im; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_11_re <= 64'sh0; // @[Cholesky_V1.scala 46:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_11_re <= io_matrixIn_11_re; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_11_im <= 64'sh0; // @[Cholesky_V1.scala 47:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_11_im <= io_matrixIn_11_im; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_12_re <= 64'sh0; // @[Cholesky_V1.scala 46:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_12_re <= io_matrixIn_12_re; // @[Cholesky_V1.scala 52:21]
    end else if (!(status <= 8'h1f)) begin // @[Cholesky_V1.scala 56:48]
      if (!(status == 8'h20)) begin // @[Cholesky_V1.scala 60:55]
        matrix_comp_reg_12_re <= _GEN_33;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_12_im <= 64'sh0; // @[Cholesky_V1.scala 47:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_12_im <= io_matrixIn_12_im; // @[Cholesky_V1.scala 52:21]
    end else if (!(status <= 8'h1f)) begin // @[Cholesky_V1.scala 56:48]
      if (!(status == 8'h20)) begin // @[Cholesky_V1.scala 60:55]
        matrix_comp_reg_12_im <= _GEN_32;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_13_re <= 64'sh0; // @[Cholesky_V1.scala 46:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_13_re <= io_matrixIn_13_re; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_13_im <= 64'sh0; // @[Cholesky_V1.scala 47:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_13_im <= io_matrixIn_13_im; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_14_re <= 64'sh0; // @[Cholesky_V1.scala 46:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_14_re <= io_matrixIn_14_re; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_14_im <= 64'sh0; // @[Cholesky_V1.scala 47:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_14_im <= io_matrixIn_14_im; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_15_re <= 64'sh0; // @[Cholesky_V1.scala 46:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_15_re <= io_matrixIn_15_re; // @[Cholesky_V1.scala 52:21]
    end
    if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      matrix_comp_reg_15_im <= 64'sh0; // @[Cholesky_V1.scala 47:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      matrix_comp_reg_15_im <= io_matrixIn_15_im; // @[Cholesky_V1.scala 52:21]
    end
    if (reset) begin // @[Cholesky_V1.scala 24:29]
      status <= 8'h0; // @[Cholesky_V1.scala 24:29]
    end else if (io_reset) begin // @[Cholesky_V1.scala 43:18]
      status <= 8'h0; // @[Cholesky_V1.scala 49:12]
    end else if (io_ready) begin // @[Cholesky_V1.scala 50:24]
      status <= 8'h1; // @[Cholesky_V1.scala 53:12]
    end else if (status <= 8'h1f) begin // @[Cholesky_V1.scala 56:48]
      status <= _status_T_1; // @[Cholesky_V1.scala 59:14]
    end else begin
      status <= _GEN_43;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  matrix_comp_reg_0_re = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  matrix_comp_reg_0_im = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  matrix_comp_reg_1_re = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  matrix_comp_reg_1_im = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  matrix_comp_reg_2_re = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  matrix_comp_reg_2_im = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  matrix_comp_reg_3_re = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  matrix_comp_reg_3_im = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  matrix_comp_reg_4_re = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  matrix_comp_reg_4_im = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  matrix_comp_reg_5_re = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  matrix_comp_reg_5_im = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  matrix_comp_reg_6_re = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  matrix_comp_reg_6_im = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  matrix_comp_reg_7_re = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  matrix_comp_reg_7_im = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  matrix_comp_reg_8_re = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  matrix_comp_reg_8_im = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  matrix_comp_reg_9_re = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  matrix_comp_reg_9_im = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  matrix_comp_reg_10_re = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  matrix_comp_reg_10_im = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  matrix_comp_reg_11_re = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  matrix_comp_reg_11_im = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  matrix_comp_reg_12_re = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  matrix_comp_reg_12_im = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  matrix_comp_reg_13_re = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  matrix_comp_reg_13_im = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  matrix_comp_reg_14_re = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  matrix_comp_reg_14_im = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  matrix_comp_reg_15_re = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  matrix_comp_reg_15_im = _RAND_31[63:0];
  _RAND_32 = {1{`RANDOM}};
  status = _RAND_32[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cholesky_v1(
  input         clock,
  input         reset,
  input         io_reset,
  input         io_ready,
  input  [63:0] io_matrixIn_0_re,
  input  [63:0] io_matrixIn_0_im,
  input  [63:0] io_matrixIn_1_re,
  input  [63:0] io_matrixIn_1_im,
  input  [63:0] io_matrixIn_2_re,
  input  [63:0] io_matrixIn_2_im,
  input  [63:0] io_matrixIn_3_re,
  input  [63:0] io_matrixIn_3_im,
  input  [63:0] io_matrixIn_4_re,
  input  [63:0] io_matrixIn_4_im,
  input  [63:0] io_matrixIn_5_re,
  input  [63:0] io_matrixIn_5_im,
  input  [63:0] io_matrixIn_6_re,
  input  [63:0] io_matrixIn_6_im,
  input  [63:0] io_matrixIn_7_re,
  input  [63:0] io_matrixIn_7_im,
  input  [63:0] io_matrixIn_8_re,
  input  [63:0] io_matrixIn_8_im,
  input  [63:0] io_matrixIn_9_re,
  input  [63:0] io_matrixIn_9_im,
  input  [63:0] io_matrixIn_10_re,
  input  [63:0] io_matrixIn_10_im,
  input  [63:0] io_matrixIn_11_re,
  input  [63:0] io_matrixIn_11_im,
  input  [63:0] io_matrixIn_12_re,
  input  [63:0] io_matrixIn_12_im,
  input  [63:0] io_matrixIn_13_re,
  input  [63:0] io_matrixIn_13_im,
  input  [63:0] io_matrixIn_14_re,
  input  [63:0] io_matrixIn_14_im,
  input  [63:0] io_matrixIn_15_re,
  input  [63:0] io_matrixIn_15_im,
  output [63:0] io_matrixOut_0_re,
  output [63:0] io_matrixOut_0_im,
  output [63:0] io_matrixOut_1_re,
  output [63:0] io_matrixOut_1_im,
  output [63:0] io_matrixOut_2_re,
  output [63:0] io_matrixOut_2_im,
  output [63:0] io_matrixOut_3_re,
  output [63:0] io_matrixOut_3_im,
  output [63:0] io_matrixOut_4_re,
  output [63:0] io_matrixOut_4_im,
  output [63:0] io_matrixOut_5_re,
  output [63:0] io_matrixOut_5_im,
  output [63:0] io_matrixOut_6_re,
  output [63:0] io_matrixOut_6_im,
  output [63:0] io_matrixOut_7_re,
  output [63:0] io_matrixOut_7_im,
  output [63:0] io_matrixOut_8_re,
  output [63:0] io_matrixOut_8_im,
  output [63:0] io_matrixOut_9_re,
  output [63:0] io_matrixOut_9_im,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  wire  cholesky_comp_unit_clock; // @[Cholesky_V1.scala 131:54]
  wire  cholesky_comp_unit_reset; // @[Cholesky_V1.scala 131:54]
  wire  cholesky_comp_unit_io_reset; // @[Cholesky_V1.scala 131:54]
  wire  cholesky_comp_unit_io_ready; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_0_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_0_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_1_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_1_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_2_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_2_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_3_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_3_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_4_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_4_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_5_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_5_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_6_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_6_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_7_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_7_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_8_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_8_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_9_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_9_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_10_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_10_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_11_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_11_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_12_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_12_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_13_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_13_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_14_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_14_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_15_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixIn_15_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_0_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_0_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_1_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_1_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_2_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_2_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_3_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_3_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_4_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_4_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_5_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_5_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_6_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_6_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_7_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_7_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_8_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_8_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_9_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_9_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_10_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_10_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_11_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_11_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_12_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_12_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_13_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_13_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_14_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_14_im; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_15_re; // @[Cholesky_V1.scala 131:54]
  wire [63:0] cholesky_comp_unit_io_matrixOut_15_im; // @[Cholesky_V1.scala 131:54]
  wire  cholesky_comp_unit_io_valid; // @[Cholesky_V1.scala 131:54]
  reg [63:0] matrix_comp_reg_0_re; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_0_im; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_1_re; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_1_im; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_2_re; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_2_im; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_3_re; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_3_im; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_4_re; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_4_im; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_5_re; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_5_im; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_6_re; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_6_im; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_7_re; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_7_im; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_8_re; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_8_im; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_9_re; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_9_im; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_10_re; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_10_im; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_11_re; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_11_im; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_12_re; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_12_im; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_13_re; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_13_im; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_14_re; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_14_im; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_15_re; // @[Cholesky_V1.scala 127:42]
  reg [63:0] matrix_comp_reg_15_im; // @[Cholesky_V1.scala 127:42]
  reg [31:0] point_index; // @[Cholesky_V1.scala 128:34]
  reg [3:0] comp_status; // @[Cholesky_V1.scala 129:34]
  wire [31:0] _T_2 = 32'h4 - point_index; // @[Cholesky_V1.scala 157:28]
  wire [32:0] _cholesky_comp_unit_io_matrixIn_0_T = {{1'd0}, point_index}; // @[Cholesky_V1.scala 158:78]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_0_T_2 = _cholesky_comp_unit_io_matrixIn_0_T[31:0] * 3'h4; // @[Cholesky_V1.scala 158:92]
  wire [34:0] _GEN_1360 = {{3'd0}, _cholesky_comp_unit_io_matrixIn_0_T[31:0]}; // @[Cholesky_V1.scala 158:98]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_0_T_6 = _cholesky_comp_unit_io_matrixIn_0_T_2 + _GEN_1360; // @[Cholesky_V1.scala 158:98]
  wire [63:0] _GEN_1 = 4'h1 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_1_im) : $signed(
    matrix_comp_reg_0_im); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_2 = 4'h2 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_2_im) : $signed(
    _GEN_1); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_3 = 4'h3 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_3_im) : $signed(
    _GEN_2); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_4 = 4'h4 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_4_im) : $signed(
    _GEN_3); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_5 = 4'h5 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_5_im) : $signed(
    _GEN_4); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_6 = 4'h6 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_6_im) : $signed(
    _GEN_5); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_7 = 4'h7 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_7_im) : $signed(
    _GEN_6); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_8 = 4'h8 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_8_im) : $signed(
    _GEN_7); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_9 = 4'h9 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_9_im) : $signed(
    _GEN_8); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_10 = 4'ha == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_10_im) : $signed(
    _GEN_9); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_11 = 4'hb == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_11_im) : $signed(
    _GEN_10); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_12 = 4'hc == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_12_im) : $signed(
    _GEN_11); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_13 = 4'hd == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_13_im) : $signed(
    _GEN_12); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_14 = 4'he == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_14_im) : $signed(
    _GEN_13); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_17 = 4'h1 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_1_re) : $signed(
    matrix_comp_reg_0_re); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_18 = 4'h2 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_2_re) : $signed(
    _GEN_17); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_19 = 4'h3 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_3_re) : $signed(
    _GEN_18); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_20 = 4'h4 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_4_re) : $signed(
    _GEN_19); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_21 = 4'h5 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_5_re) : $signed(
    _GEN_20); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_22 = 4'h6 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_6_re) : $signed(
    _GEN_21); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_23 = 4'h7 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_7_re) : $signed(
    _GEN_22); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_24 = 4'h8 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_8_re) : $signed(
    _GEN_23); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_25 = 4'h9 == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_9_re) : $signed(
    _GEN_24); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_26 = 4'ha == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_10_re) : $signed(
    _GEN_25); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_27 = 4'hb == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_11_re) : $signed(
    _GEN_26); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_28 = 4'hc == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_12_re) : $signed(
    _GEN_27); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_29 = 4'hd == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_13_re) : $signed(
    _GEN_28); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_30 = 4'he == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_14_re) : $signed(
    _GEN_29); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_31 = 4'hf == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(matrix_comp_reg_15_re) : $signed(
    _GEN_30); // @[Cholesky_V1.scala 158:{55,55}]
  wire [31:0] _cholesky_comp_unit_io_matrixIn_1_T_4 = 32'h1 + point_index; // @[Cholesky_V1.scala 158:104]
  wire [34:0] _GEN_1361 = {{3'd0}, _cholesky_comp_unit_io_matrixIn_1_T_4}; // @[Cholesky_V1.scala 158:98]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_1_T_6 = _cholesky_comp_unit_io_matrixIn_0_T_2 + _GEN_1361; // @[Cholesky_V1.scala 158:98]
  wire [63:0] _GEN_35 = 4'h1 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_1_im) : $signed(
    matrix_comp_reg_0_im); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_36 = 4'h2 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_2_im) : $signed(
    _GEN_35); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_37 = 4'h3 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_3_im) : $signed(
    _GEN_36); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_38 = 4'h4 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_4_im) : $signed(
    _GEN_37); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_39 = 4'h5 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_5_im) : $signed(
    _GEN_38); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_40 = 4'h6 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_6_im) : $signed(
    _GEN_39); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_41 = 4'h7 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_7_im) : $signed(
    _GEN_40); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_42 = 4'h8 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_8_im) : $signed(
    _GEN_41); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_43 = 4'h9 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_9_im) : $signed(
    _GEN_42); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_44 = 4'ha == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_10_im) : $signed(
    _GEN_43); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_45 = 4'hb == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_11_im) : $signed(
    _GEN_44); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_46 = 4'hc == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_12_im) : $signed(
    _GEN_45); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_47 = 4'hd == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_13_im) : $signed(
    _GEN_46); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_48 = 4'he == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_14_im) : $signed(
    _GEN_47); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_51 = 4'h1 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_1_re) : $signed(
    matrix_comp_reg_0_re); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_52 = 4'h2 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_2_re) : $signed(
    _GEN_51); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_53 = 4'h3 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_3_re) : $signed(
    _GEN_52); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_54 = 4'h4 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_4_re) : $signed(
    _GEN_53); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_55 = 4'h5 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_5_re) : $signed(
    _GEN_54); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_56 = 4'h6 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_6_re) : $signed(
    _GEN_55); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_57 = 4'h7 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_7_re) : $signed(
    _GEN_56); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_58 = 4'h8 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_8_re) : $signed(
    _GEN_57); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_59 = 4'h9 == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_9_re) : $signed(
    _GEN_58); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_60 = 4'ha == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_10_re) : $signed(
    _GEN_59); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_61 = 4'hb == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_11_re) : $signed(
    _GEN_60); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_62 = 4'hc == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_12_re) : $signed(
    _GEN_61); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_63 = 4'hd == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_13_re) : $signed(
    _GEN_62); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_64 = 4'he == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_14_re) : $signed(
    _GEN_63); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_65 = 4'hf == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(matrix_comp_reg_15_re) : $signed(
    _GEN_64); // @[Cholesky_V1.scala 158:{55,55}]
  wire [31:0] _cholesky_comp_unit_io_matrixIn_2_T_4 = 32'h2 + point_index; // @[Cholesky_V1.scala 158:104]
  wire [34:0] _GEN_1362 = {{3'd0}, _cholesky_comp_unit_io_matrixIn_2_T_4}; // @[Cholesky_V1.scala 158:98]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_2_T_6 = _cholesky_comp_unit_io_matrixIn_0_T_2 + _GEN_1362; // @[Cholesky_V1.scala 158:98]
  wire [63:0] _GEN_69 = 4'h1 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_1_im) : $signed(
    matrix_comp_reg_0_im); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_70 = 4'h2 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_2_im) : $signed(
    _GEN_69); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_71 = 4'h3 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_3_im) : $signed(
    _GEN_70); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_72 = 4'h4 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_4_im) : $signed(
    _GEN_71); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_73 = 4'h5 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_5_im) : $signed(
    _GEN_72); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_74 = 4'h6 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_6_im) : $signed(
    _GEN_73); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_75 = 4'h7 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_7_im) : $signed(
    _GEN_74); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_76 = 4'h8 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_8_im) : $signed(
    _GEN_75); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_77 = 4'h9 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_9_im) : $signed(
    _GEN_76); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_78 = 4'ha == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_10_im) : $signed(
    _GEN_77); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_79 = 4'hb == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_11_im) : $signed(
    _GEN_78); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_80 = 4'hc == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_12_im) : $signed(
    _GEN_79); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_81 = 4'hd == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_13_im) : $signed(
    _GEN_80); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_82 = 4'he == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_14_im) : $signed(
    _GEN_81); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_85 = 4'h1 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_1_re) : $signed(
    matrix_comp_reg_0_re); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_86 = 4'h2 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_2_re) : $signed(
    _GEN_85); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_87 = 4'h3 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_3_re) : $signed(
    _GEN_86); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_88 = 4'h4 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_4_re) : $signed(
    _GEN_87); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_89 = 4'h5 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_5_re) : $signed(
    _GEN_88); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_90 = 4'h6 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_6_re) : $signed(
    _GEN_89); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_91 = 4'h7 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_7_re) : $signed(
    _GEN_90); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_92 = 4'h8 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_8_re) : $signed(
    _GEN_91); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_93 = 4'h9 == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_9_re) : $signed(
    _GEN_92); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_94 = 4'ha == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_10_re) : $signed(
    _GEN_93); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_95 = 4'hb == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_11_re) : $signed(
    _GEN_94); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_96 = 4'hc == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_12_re) : $signed(
    _GEN_95); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_97 = 4'hd == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_13_re) : $signed(
    _GEN_96); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_98 = 4'he == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_14_re) : $signed(
    _GEN_97); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_99 = 4'hf == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(matrix_comp_reg_15_re) : $signed(
    _GEN_98); // @[Cholesky_V1.scala 158:{55,55}]
  wire [31:0] _cholesky_comp_unit_io_matrixIn_3_T_4 = 32'h3 + point_index; // @[Cholesky_V1.scala 158:104]
  wire [34:0] _GEN_1363 = {{3'd0}, _cholesky_comp_unit_io_matrixIn_3_T_4}; // @[Cholesky_V1.scala 158:98]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_3_T_6 = _cholesky_comp_unit_io_matrixIn_0_T_2 + _GEN_1363; // @[Cholesky_V1.scala 158:98]
  wire [63:0] _GEN_103 = 4'h1 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_1_im) : $signed(
    matrix_comp_reg_0_im); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_104 = 4'h2 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_2_im) : $signed(
    _GEN_103); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_105 = 4'h3 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_3_im) : $signed(
    _GEN_104); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_106 = 4'h4 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_4_im) : $signed(
    _GEN_105); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_107 = 4'h5 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_5_im) : $signed(
    _GEN_106); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_108 = 4'h6 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_6_im) : $signed(
    _GEN_107); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_109 = 4'h7 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_7_im) : $signed(
    _GEN_108); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_110 = 4'h8 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_8_im) : $signed(
    _GEN_109); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_111 = 4'h9 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_9_im) : $signed(
    _GEN_110); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_112 = 4'ha == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_10_im) : $signed(
    _GEN_111); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_113 = 4'hb == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_11_im) : $signed(
    _GEN_112); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_114 = 4'hc == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_12_im) : $signed(
    _GEN_113); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_115 = 4'hd == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_13_im) : $signed(
    _GEN_114); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_116 = 4'he == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_14_im) : $signed(
    _GEN_115); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_119 = 4'h1 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_1_re) : $signed(
    matrix_comp_reg_0_re); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_120 = 4'h2 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_2_re) : $signed(
    _GEN_119); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_121 = 4'h3 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_3_re) : $signed(
    _GEN_120); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_122 = 4'h4 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_4_re) : $signed(
    _GEN_121); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_123 = 4'h5 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_5_re) : $signed(
    _GEN_122); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_124 = 4'h6 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_6_re) : $signed(
    _GEN_123); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_125 = 4'h7 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_7_re) : $signed(
    _GEN_124); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_126 = 4'h8 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_8_re) : $signed(
    _GEN_125); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_127 = 4'h9 == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_9_re) : $signed(
    _GEN_126); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_128 = 4'ha == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_10_re) : $signed(
    _GEN_127); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_129 = 4'hb == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_11_re) : $signed(
    _GEN_128); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_130 = 4'hc == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_12_re) : $signed(
    _GEN_129); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_131 = 4'hd == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_13_re) : $signed(
    _GEN_130); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_132 = 4'he == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_14_re) : $signed(
    _GEN_131); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_133 = 4'hf == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(matrix_comp_reg_15_re) : $signed(
    _GEN_132); // @[Cholesky_V1.scala 158:{55,55}]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_4_T_2 = _cholesky_comp_unit_io_matrixIn_1_T_4 * 3'h4; // @[Cholesky_V1.scala 158:92]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_4_T_6 = _cholesky_comp_unit_io_matrixIn_4_T_2 + _GEN_1360; // @[Cholesky_V1.scala 158:98]
  wire [63:0] _GEN_137 = 4'h1 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_1_im) : $signed(
    matrix_comp_reg_0_im); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_138 = 4'h2 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_2_im) : $signed(
    _GEN_137); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_139 = 4'h3 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_3_im) : $signed(
    _GEN_138); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_140 = 4'h4 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_4_im) : $signed(
    _GEN_139); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_141 = 4'h5 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_5_im) : $signed(
    _GEN_140); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_142 = 4'h6 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_6_im) : $signed(
    _GEN_141); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_143 = 4'h7 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_7_im) : $signed(
    _GEN_142); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_144 = 4'h8 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_8_im) : $signed(
    _GEN_143); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_145 = 4'h9 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_9_im) : $signed(
    _GEN_144); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_146 = 4'ha == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_10_im) : $signed(
    _GEN_145); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_147 = 4'hb == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_11_im) : $signed(
    _GEN_146); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_148 = 4'hc == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_12_im) : $signed(
    _GEN_147); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_149 = 4'hd == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_13_im) : $signed(
    _GEN_148); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_150 = 4'he == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_14_im) : $signed(
    _GEN_149); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_153 = 4'h1 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_1_re) : $signed(
    matrix_comp_reg_0_re); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_154 = 4'h2 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_2_re) : $signed(
    _GEN_153); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_155 = 4'h3 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_3_re) : $signed(
    _GEN_154); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_156 = 4'h4 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_4_re) : $signed(
    _GEN_155); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_157 = 4'h5 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_5_re) : $signed(
    _GEN_156); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_158 = 4'h6 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_6_re) : $signed(
    _GEN_157); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_159 = 4'h7 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_7_re) : $signed(
    _GEN_158); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_160 = 4'h8 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_8_re) : $signed(
    _GEN_159); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_161 = 4'h9 == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_9_re) : $signed(
    _GEN_160); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_162 = 4'ha == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_10_re) : $signed(
    _GEN_161); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_163 = 4'hb == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_11_re) : $signed(
    _GEN_162); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_164 = 4'hc == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_12_re) : $signed(
    _GEN_163); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_165 = 4'hd == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_13_re) : $signed(
    _GEN_164); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_166 = 4'he == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_14_re) : $signed(
    _GEN_165); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_167 = 4'hf == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(matrix_comp_reg_15_re) : $signed(
    _GEN_166); // @[Cholesky_V1.scala 158:{55,55}]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_5_T_6 = _cholesky_comp_unit_io_matrixIn_4_T_2 + _GEN_1361; // @[Cholesky_V1.scala 158:98]
  wire [63:0] _GEN_171 = 4'h1 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_1_im) : $signed(
    matrix_comp_reg_0_im); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_172 = 4'h2 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_2_im) : $signed(
    _GEN_171); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_173 = 4'h3 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_3_im) : $signed(
    _GEN_172); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_174 = 4'h4 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_4_im) : $signed(
    _GEN_173); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_175 = 4'h5 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_5_im) : $signed(
    _GEN_174); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_176 = 4'h6 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_6_im) : $signed(
    _GEN_175); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_177 = 4'h7 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_7_im) : $signed(
    _GEN_176); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_178 = 4'h8 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_8_im) : $signed(
    _GEN_177); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_179 = 4'h9 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_9_im) : $signed(
    _GEN_178); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_180 = 4'ha == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_10_im) : $signed(
    _GEN_179); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_181 = 4'hb == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_11_im) : $signed(
    _GEN_180); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_182 = 4'hc == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_12_im) : $signed(
    _GEN_181); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_183 = 4'hd == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_13_im) : $signed(
    _GEN_182); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_184 = 4'he == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_14_im) : $signed(
    _GEN_183); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_187 = 4'h1 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_1_re) : $signed(
    matrix_comp_reg_0_re); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_188 = 4'h2 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_2_re) : $signed(
    _GEN_187); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_189 = 4'h3 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_3_re) : $signed(
    _GEN_188); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_190 = 4'h4 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_4_re) : $signed(
    _GEN_189); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_191 = 4'h5 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_5_re) : $signed(
    _GEN_190); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_192 = 4'h6 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_6_re) : $signed(
    _GEN_191); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_193 = 4'h7 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_7_re) : $signed(
    _GEN_192); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_194 = 4'h8 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_8_re) : $signed(
    _GEN_193); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_195 = 4'h9 == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_9_re) : $signed(
    _GEN_194); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_196 = 4'ha == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_10_re) : $signed(
    _GEN_195); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_197 = 4'hb == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_11_re) : $signed(
    _GEN_196); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_198 = 4'hc == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_12_re) : $signed(
    _GEN_197); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_199 = 4'hd == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_13_re) : $signed(
    _GEN_198); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_200 = 4'he == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_14_re) : $signed(
    _GEN_199); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_201 = 4'hf == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(matrix_comp_reg_15_re) : $signed(
    _GEN_200); // @[Cholesky_V1.scala 158:{55,55}]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_6_T_6 = _cholesky_comp_unit_io_matrixIn_4_T_2 + _GEN_1362; // @[Cholesky_V1.scala 158:98]
  wire [63:0] _GEN_205 = 4'h1 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_1_im) : $signed(
    matrix_comp_reg_0_im); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_206 = 4'h2 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_2_im) : $signed(
    _GEN_205); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_207 = 4'h3 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_3_im) : $signed(
    _GEN_206); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_208 = 4'h4 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_4_im) : $signed(
    _GEN_207); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_209 = 4'h5 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_5_im) : $signed(
    _GEN_208); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_210 = 4'h6 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_6_im) : $signed(
    _GEN_209); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_211 = 4'h7 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_7_im) : $signed(
    _GEN_210); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_212 = 4'h8 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_8_im) : $signed(
    _GEN_211); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_213 = 4'h9 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_9_im) : $signed(
    _GEN_212); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_214 = 4'ha == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_10_im) : $signed(
    _GEN_213); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_215 = 4'hb == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_11_im) : $signed(
    _GEN_214); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_216 = 4'hc == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_12_im) : $signed(
    _GEN_215); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_217 = 4'hd == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_13_im) : $signed(
    _GEN_216); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_218 = 4'he == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_14_im) : $signed(
    _GEN_217); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_221 = 4'h1 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_1_re) : $signed(
    matrix_comp_reg_0_re); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_222 = 4'h2 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_2_re) : $signed(
    _GEN_221); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_223 = 4'h3 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_3_re) : $signed(
    _GEN_222); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_224 = 4'h4 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_4_re) : $signed(
    _GEN_223); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_225 = 4'h5 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_5_re) : $signed(
    _GEN_224); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_226 = 4'h6 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_6_re) : $signed(
    _GEN_225); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_227 = 4'h7 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_7_re) : $signed(
    _GEN_226); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_228 = 4'h8 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_8_re) : $signed(
    _GEN_227); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_229 = 4'h9 == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_9_re) : $signed(
    _GEN_228); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_230 = 4'ha == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_10_re) : $signed(
    _GEN_229); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_231 = 4'hb == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_11_re) : $signed(
    _GEN_230); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_232 = 4'hc == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_12_re) : $signed(
    _GEN_231); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_233 = 4'hd == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_13_re) : $signed(
    _GEN_232); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_234 = 4'he == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_14_re) : $signed(
    _GEN_233); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_235 = 4'hf == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(matrix_comp_reg_15_re) : $signed(
    _GEN_234); // @[Cholesky_V1.scala 158:{55,55}]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_7_T_6 = _cholesky_comp_unit_io_matrixIn_4_T_2 + _GEN_1363; // @[Cholesky_V1.scala 158:98]
  wire [63:0] _GEN_239 = 4'h1 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_1_im) : $signed(
    matrix_comp_reg_0_im); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_240 = 4'h2 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_2_im) : $signed(
    _GEN_239); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_241 = 4'h3 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_3_im) : $signed(
    _GEN_240); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_242 = 4'h4 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_4_im) : $signed(
    _GEN_241); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_243 = 4'h5 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_5_im) : $signed(
    _GEN_242); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_244 = 4'h6 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_6_im) : $signed(
    _GEN_243); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_245 = 4'h7 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_7_im) : $signed(
    _GEN_244); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_246 = 4'h8 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_8_im) : $signed(
    _GEN_245); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_247 = 4'h9 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_9_im) : $signed(
    _GEN_246); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_248 = 4'ha == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_10_im) : $signed(
    _GEN_247); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_249 = 4'hb == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_11_im) : $signed(
    _GEN_248); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_250 = 4'hc == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_12_im) : $signed(
    _GEN_249); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_251 = 4'hd == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_13_im) : $signed(
    _GEN_250); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_252 = 4'he == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_14_im) : $signed(
    _GEN_251); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_255 = 4'h1 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_1_re) : $signed(
    matrix_comp_reg_0_re); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_256 = 4'h2 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_2_re) : $signed(
    _GEN_255); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_257 = 4'h3 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_3_re) : $signed(
    _GEN_256); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_258 = 4'h4 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_4_re) : $signed(
    _GEN_257); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_259 = 4'h5 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_5_re) : $signed(
    _GEN_258); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_260 = 4'h6 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_6_re) : $signed(
    _GEN_259); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_261 = 4'h7 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_7_re) : $signed(
    _GEN_260); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_262 = 4'h8 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_8_re) : $signed(
    _GEN_261); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_263 = 4'h9 == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_9_re) : $signed(
    _GEN_262); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_264 = 4'ha == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_10_re) : $signed(
    _GEN_263); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_265 = 4'hb == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_11_re) : $signed(
    _GEN_264); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_266 = 4'hc == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_12_re) : $signed(
    _GEN_265); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_267 = 4'hd == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_13_re) : $signed(
    _GEN_266); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_268 = 4'he == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_14_re) : $signed(
    _GEN_267); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_269 = 4'hf == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(matrix_comp_reg_15_re) : $signed(
    _GEN_268); // @[Cholesky_V1.scala 158:{55,55}]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_8_T_2 = _cholesky_comp_unit_io_matrixIn_2_T_4 * 3'h4; // @[Cholesky_V1.scala 158:92]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_8_T_6 = _cholesky_comp_unit_io_matrixIn_8_T_2 + _GEN_1360; // @[Cholesky_V1.scala 158:98]
  wire [63:0] _GEN_273 = 4'h1 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_1_im) : $signed(
    matrix_comp_reg_0_im); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_274 = 4'h2 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_2_im) : $signed(
    _GEN_273); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_275 = 4'h3 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_3_im) : $signed(
    _GEN_274); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_276 = 4'h4 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_4_im) : $signed(
    _GEN_275); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_277 = 4'h5 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_5_im) : $signed(
    _GEN_276); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_278 = 4'h6 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_6_im) : $signed(
    _GEN_277); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_279 = 4'h7 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_7_im) : $signed(
    _GEN_278); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_280 = 4'h8 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_8_im) : $signed(
    _GEN_279); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_281 = 4'h9 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_9_im) : $signed(
    _GEN_280); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_282 = 4'ha == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_10_im) : $signed(
    _GEN_281); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_283 = 4'hb == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_11_im) : $signed(
    _GEN_282); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_284 = 4'hc == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_12_im) : $signed(
    _GEN_283); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_285 = 4'hd == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_13_im) : $signed(
    _GEN_284); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_286 = 4'he == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_14_im) : $signed(
    _GEN_285); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_289 = 4'h1 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_1_re) : $signed(
    matrix_comp_reg_0_re); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_290 = 4'h2 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_2_re) : $signed(
    _GEN_289); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_291 = 4'h3 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_3_re) : $signed(
    _GEN_290); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_292 = 4'h4 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_4_re) : $signed(
    _GEN_291); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_293 = 4'h5 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_5_re) : $signed(
    _GEN_292); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_294 = 4'h6 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_6_re) : $signed(
    _GEN_293); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_295 = 4'h7 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_7_re) : $signed(
    _GEN_294); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_296 = 4'h8 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_8_re) : $signed(
    _GEN_295); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_297 = 4'h9 == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_9_re) : $signed(
    _GEN_296); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_298 = 4'ha == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_10_re) : $signed(
    _GEN_297); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_299 = 4'hb == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_11_re) : $signed(
    _GEN_298); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_300 = 4'hc == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_12_re) : $signed(
    _GEN_299); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_301 = 4'hd == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_13_re) : $signed(
    _GEN_300); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_302 = 4'he == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_14_re) : $signed(
    _GEN_301); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_303 = 4'hf == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(matrix_comp_reg_15_re) : $signed(
    _GEN_302); // @[Cholesky_V1.scala 158:{55,55}]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_9_T_6 = _cholesky_comp_unit_io_matrixIn_8_T_2 + _GEN_1361; // @[Cholesky_V1.scala 158:98]
  wire [63:0] _GEN_307 = 4'h1 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_1_im) : $signed(
    matrix_comp_reg_0_im); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_308 = 4'h2 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_2_im) : $signed(
    _GEN_307); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_309 = 4'h3 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_3_im) : $signed(
    _GEN_308); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_310 = 4'h4 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_4_im) : $signed(
    _GEN_309); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_311 = 4'h5 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_5_im) : $signed(
    _GEN_310); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_312 = 4'h6 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_6_im) : $signed(
    _GEN_311); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_313 = 4'h7 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_7_im) : $signed(
    _GEN_312); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_314 = 4'h8 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_8_im) : $signed(
    _GEN_313); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_315 = 4'h9 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_9_im) : $signed(
    _GEN_314); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_316 = 4'ha == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_10_im) : $signed(
    _GEN_315); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_317 = 4'hb == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_11_im) : $signed(
    _GEN_316); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_318 = 4'hc == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_12_im) : $signed(
    _GEN_317); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_319 = 4'hd == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_13_im) : $signed(
    _GEN_318); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_320 = 4'he == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_14_im) : $signed(
    _GEN_319); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_323 = 4'h1 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_1_re) : $signed(
    matrix_comp_reg_0_re); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_324 = 4'h2 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_2_re) : $signed(
    _GEN_323); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_325 = 4'h3 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_3_re) : $signed(
    _GEN_324); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_326 = 4'h4 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_4_re) : $signed(
    _GEN_325); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_327 = 4'h5 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_5_re) : $signed(
    _GEN_326); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_328 = 4'h6 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_6_re) : $signed(
    _GEN_327); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_329 = 4'h7 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_7_re) : $signed(
    _GEN_328); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_330 = 4'h8 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_8_re) : $signed(
    _GEN_329); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_331 = 4'h9 == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_9_re) : $signed(
    _GEN_330); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_332 = 4'ha == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_10_re) : $signed(
    _GEN_331); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_333 = 4'hb == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_11_re) : $signed(
    _GEN_332); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_334 = 4'hc == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_12_re) : $signed(
    _GEN_333); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_335 = 4'hd == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_13_re) : $signed(
    _GEN_334); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_336 = 4'he == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_14_re) : $signed(
    _GEN_335); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_337 = 4'hf == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(matrix_comp_reg_15_re) : $signed(
    _GEN_336); // @[Cholesky_V1.scala 158:{55,55}]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_10_T_6 = _cholesky_comp_unit_io_matrixIn_8_T_2 + _GEN_1362; // @[Cholesky_V1.scala 158:98]
  wire [63:0] _GEN_341 = 4'h1 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_1_im) : $signed(
    matrix_comp_reg_0_im); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_342 = 4'h2 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_2_im) : $signed(
    _GEN_341); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_343 = 4'h3 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_3_im) : $signed(
    _GEN_342); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_344 = 4'h4 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_4_im) : $signed(
    _GEN_343); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_345 = 4'h5 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_5_im) : $signed(
    _GEN_344); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_346 = 4'h6 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_6_im) : $signed(
    _GEN_345); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_347 = 4'h7 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_7_im) : $signed(
    _GEN_346); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_348 = 4'h8 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_8_im) : $signed(
    _GEN_347); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_349 = 4'h9 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_9_im) : $signed(
    _GEN_348); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_350 = 4'ha == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_10_im) : $signed(
    _GEN_349); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_351 = 4'hb == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_11_im) : $signed(
    _GEN_350); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_352 = 4'hc == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_12_im) : $signed(
    _GEN_351); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_353 = 4'hd == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_13_im) : $signed(
    _GEN_352); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_354 = 4'he == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_14_im) : $signed(
    _GEN_353); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_357 = 4'h1 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_1_re) : $signed(
    matrix_comp_reg_0_re); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_358 = 4'h2 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_2_re) : $signed(
    _GEN_357); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_359 = 4'h3 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_3_re) : $signed(
    _GEN_358); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_360 = 4'h4 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_4_re) : $signed(
    _GEN_359); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_361 = 4'h5 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_5_re) : $signed(
    _GEN_360); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_362 = 4'h6 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_6_re) : $signed(
    _GEN_361); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_363 = 4'h7 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_7_re) : $signed(
    _GEN_362); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_364 = 4'h8 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_8_re) : $signed(
    _GEN_363); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_365 = 4'h9 == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_9_re) : $signed(
    _GEN_364); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_366 = 4'ha == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_10_re) : $signed(
    _GEN_365); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_367 = 4'hb == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_11_re) : $signed(
    _GEN_366); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_368 = 4'hc == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_12_re) : $signed(
    _GEN_367); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_369 = 4'hd == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_13_re) : $signed(
    _GEN_368); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_370 = 4'he == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_14_re) : $signed(
    _GEN_369); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_371 = 4'hf == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(matrix_comp_reg_15_re) : $signed(
    _GEN_370); // @[Cholesky_V1.scala 158:{55,55}]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_11_T_6 = _cholesky_comp_unit_io_matrixIn_8_T_2 + _GEN_1363; // @[Cholesky_V1.scala 158:98]
  wire [63:0] _GEN_375 = 4'h1 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_1_im) : $signed(
    matrix_comp_reg_0_im); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_376 = 4'h2 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_2_im) : $signed(
    _GEN_375); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_377 = 4'h3 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_3_im) : $signed(
    _GEN_376); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_378 = 4'h4 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_4_im) : $signed(
    _GEN_377); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_379 = 4'h5 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_5_im) : $signed(
    _GEN_378); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_380 = 4'h6 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_6_im) : $signed(
    _GEN_379); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_381 = 4'h7 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_7_im) : $signed(
    _GEN_380); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_382 = 4'h8 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_8_im) : $signed(
    _GEN_381); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_383 = 4'h9 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_9_im) : $signed(
    _GEN_382); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_384 = 4'ha == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_10_im) : $signed(
    _GEN_383); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_385 = 4'hb == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_11_im) : $signed(
    _GEN_384); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_386 = 4'hc == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_12_im) : $signed(
    _GEN_385); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_387 = 4'hd == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_13_im) : $signed(
    _GEN_386); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_388 = 4'he == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_14_im) : $signed(
    _GEN_387); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_391 = 4'h1 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_1_re) : $signed(
    matrix_comp_reg_0_re); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_392 = 4'h2 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_2_re) : $signed(
    _GEN_391); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_393 = 4'h3 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_3_re) : $signed(
    _GEN_392); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_394 = 4'h4 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_4_re) : $signed(
    _GEN_393); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_395 = 4'h5 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_5_re) : $signed(
    _GEN_394); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_396 = 4'h6 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_6_re) : $signed(
    _GEN_395); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_397 = 4'h7 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_7_re) : $signed(
    _GEN_396); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_398 = 4'h8 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_8_re) : $signed(
    _GEN_397); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_399 = 4'h9 == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_9_re) : $signed(
    _GEN_398); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_400 = 4'ha == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_10_re) : $signed(
    _GEN_399); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_401 = 4'hb == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_11_re) : $signed(
    _GEN_400); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_402 = 4'hc == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_12_re) : $signed(
    _GEN_401); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_403 = 4'hd == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_13_re) : $signed(
    _GEN_402); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_404 = 4'he == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_14_re) : $signed(
    _GEN_403); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_405 = 4'hf == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(matrix_comp_reg_15_re) : $signed(
    _GEN_404); // @[Cholesky_V1.scala 158:{55,55}]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_12_T_2 = _cholesky_comp_unit_io_matrixIn_3_T_4 * 3'h4; // @[Cholesky_V1.scala 158:92]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_12_T_6 = _cholesky_comp_unit_io_matrixIn_12_T_2 + _GEN_1360; // @[Cholesky_V1.scala 158:98]
  wire [63:0] _GEN_409 = 4'h1 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_1_im) : $signed(
    matrix_comp_reg_0_im); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_410 = 4'h2 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_2_im) : $signed(
    _GEN_409); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_411 = 4'h3 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_3_im) : $signed(
    _GEN_410); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_412 = 4'h4 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_4_im) : $signed(
    _GEN_411); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_413 = 4'h5 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_5_im) : $signed(
    _GEN_412); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_414 = 4'h6 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_6_im) : $signed(
    _GEN_413); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_415 = 4'h7 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_7_im) : $signed(
    _GEN_414); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_416 = 4'h8 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_8_im) : $signed(
    _GEN_415); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_417 = 4'h9 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_9_im) : $signed(
    _GEN_416); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_418 = 4'ha == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_10_im) : $signed(
    _GEN_417); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_419 = 4'hb == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_11_im) : $signed(
    _GEN_418); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_420 = 4'hc == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_12_im) : $signed(
    _GEN_419); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_421 = 4'hd == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_13_im) : $signed(
    _GEN_420); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_422 = 4'he == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_14_im) : $signed(
    _GEN_421); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_425 = 4'h1 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_1_re) : $signed(
    matrix_comp_reg_0_re); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_426 = 4'h2 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_2_re) : $signed(
    _GEN_425); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_427 = 4'h3 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_3_re) : $signed(
    _GEN_426); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_428 = 4'h4 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_4_re) : $signed(
    _GEN_427); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_429 = 4'h5 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_5_re) : $signed(
    _GEN_428); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_430 = 4'h6 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_6_re) : $signed(
    _GEN_429); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_431 = 4'h7 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_7_re) : $signed(
    _GEN_430); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_432 = 4'h8 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_8_re) : $signed(
    _GEN_431); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_433 = 4'h9 == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_9_re) : $signed(
    _GEN_432); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_434 = 4'ha == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_10_re) : $signed(
    _GEN_433); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_435 = 4'hb == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_11_re) : $signed(
    _GEN_434); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_436 = 4'hc == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_12_re) : $signed(
    _GEN_435); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_437 = 4'hd == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_13_re) : $signed(
    _GEN_436); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_438 = 4'he == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_14_re) : $signed(
    _GEN_437); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_439 = 4'hf == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(matrix_comp_reg_15_re) : $signed(
    _GEN_438); // @[Cholesky_V1.scala 158:{55,55}]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_13_T_6 = _cholesky_comp_unit_io_matrixIn_12_T_2 + _GEN_1361; // @[Cholesky_V1.scala 158:98]
  wire [63:0] _GEN_443 = 4'h1 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_1_im) : $signed(
    matrix_comp_reg_0_im); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_444 = 4'h2 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_2_im) : $signed(
    _GEN_443); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_445 = 4'h3 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_3_im) : $signed(
    _GEN_444); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_446 = 4'h4 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_4_im) : $signed(
    _GEN_445); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_447 = 4'h5 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_5_im) : $signed(
    _GEN_446); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_448 = 4'h6 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_6_im) : $signed(
    _GEN_447); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_449 = 4'h7 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_7_im) : $signed(
    _GEN_448); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_450 = 4'h8 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_8_im) : $signed(
    _GEN_449); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_451 = 4'h9 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_9_im) : $signed(
    _GEN_450); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_452 = 4'ha == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_10_im) : $signed(
    _GEN_451); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_453 = 4'hb == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_11_im) : $signed(
    _GEN_452); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_454 = 4'hc == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_12_im) : $signed(
    _GEN_453); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_455 = 4'hd == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_13_im) : $signed(
    _GEN_454); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_456 = 4'he == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_14_im) : $signed(
    _GEN_455); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_459 = 4'h1 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_1_re) : $signed(
    matrix_comp_reg_0_re); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_460 = 4'h2 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_2_re) : $signed(
    _GEN_459); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_461 = 4'h3 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_3_re) : $signed(
    _GEN_460); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_462 = 4'h4 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_4_re) : $signed(
    _GEN_461); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_463 = 4'h5 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_5_re) : $signed(
    _GEN_462); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_464 = 4'h6 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_6_re) : $signed(
    _GEN_463); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_465 = 4'h7 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_7_re) : $signed(
    _GEN_464); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_466 = 4'h8 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_8_re) : $signed(
    _GEN_465); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_467 = 4'h9 == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_9_re) : $signed(
    _GEN_466); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_468 = 4'ha == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_10_re) : $signed(
    _GEN_467); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_469 = 4'hb == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_11_re) : $signed(
    _GEN_468); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_470 = 4'hc == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_12_re) : $signed(
    _GEN_469); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_471 = 4'hd == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_13_re) : $signed(
    _GEN_470); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_472 = 4'he == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_14_re) : $signed(
    _GEN_471); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_473 = 4'hf == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(matrix_comp_reg_15_re) : $signed(
    _GEN_472); // @[Cholesky_V1.scala 158:{55,55}]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_14_T_6 = _cholesky_comp_unit_io_matrixIn_12_T_2 + _GEN_1362; // @[Cholesky_V1.scala 158:98]
  wire [63:0] _GEN_477 = 4'h1 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_1_im) : $signed(
    matrix_comp_reg_0_im); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_478 = 4'h2 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_2_im) : $signed(
    _GEN_477); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_479 = 4'h3 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_3_im) : $signed(
    _GEN_478); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_480 = 4'h4 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_4_im) : $signed(
    _GEN_479); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_481 = 4'h5 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_5_im) : $signed(
    _GEN_480); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_482 = 4'h6 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_6_im) : $signed(
    _GEN_481); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_483 = 4'h7 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_7_im) : $signed(
    _GEN_482); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_484 = 4'h8 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_8_im) : $signed(
    _GEN_483); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_485 = 4'h9 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_9_im) : $signed(
    _GEN_484); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_486 = 4'ha == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_10_im) : $signed(
    _GEN_485); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_487 = 4'hb == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_11_im) : $signed(
    _GEN_486); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_488 = 4'hc == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_12_im) : $signed(
    _GEN_487); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_489 = 4'hd == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_13_im) : $signed(
    _GEN_488); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_490 = 4'he == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_14_im) : $signed(
    _GEN_489); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_493 = 4'h1 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_1_re) : $signed(
    matrix_comp_reg_0_re); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_494 = 4'h2 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_2_re) : $signed(
    _GEN_493); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_495 = 4'h3 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_3_re) : $signed(
    _GEN_494); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_496 = 4'h4 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_4_re) : $signed(
    _GEN_495); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_497 = 4'h5 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_5_re) : $signed(
    _GEN_496); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_498 = 4'h6 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_6_re) : $signed(
    _GEN_497); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_499 = 4'h7 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_7_re) : $signed(
    _GEN_498); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_500 = 4'h8 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_8_re) : $signed(
    _GEN_499); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_501 = 4'h9 == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_9_re) : $signed(
    _GEN_500); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_502 = 4'ha == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_10_re) : $signed(
    _GEN_501); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_503 = 4'hb == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_11_re) : $signed(
    _GEN_502); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_504 = 4'hc == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_12_re) : $signed(
    _GEN_503); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_505 = 4'hd == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_13_re) : $signed(
    _GEN_504); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_506 = 4'he == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_14_re) : $signed(
    _GEN_505); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_507 = 4'hf == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(matrix_comp_reg_15_re) : $signed(
    _GEN_506); // @[Cholesky_V1.scala 158:{55,55}]
  wire [34:0] _cholesky_comp_unit_io_matrixIn_15_T_6 = _cholesky_comp_unit_io_matrixIn_12_T_2 + _GEN_1363; // @[Cholesky_V1.scala 158:98]
  wire [63:0] _GEN_511 = 4'h1 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_1_im) : $signed(
    matrix_comp_reg_0_im); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_512 = 4'h2 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_2_im) : $signed(
    _GEN_511); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_513 = 4'h3 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_3_im) : $signed(
    _GEN_512); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_514 = 4'h4 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_4_im) : $signed(
    _GEN_513); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_515 = 4'h5 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_5_im) : $signed(
    _GEN_514); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_516 = 4'h6 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_6_im) : $signed(
    _GEN_515); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_517 = 4'h7 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_7_im) : $signed(
    _GEN_516); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_518 = 4'h8 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_8_im) : $signed(
    _GEN_517); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_519 = 4'h9 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_9_im) : $signed(
    _GEN_518); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_520 = 4'ha == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_10_im) : $signed(
    _GEN_519); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_521 = 4'hb == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_11_im) : $signed(
    _GEN_520); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_522 = 4'hc == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_12_im) : $signed(
    _GEN_521); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_523 = 4'hd == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_13_im) : $signed(
    _GEN_522); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_524 = 4'he == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_14_im) : $signed(
    _GEN_523); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_527 = 4'h1 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_1_re) : $signed(
    matrix_comp_reg_0_re); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_528 = 4'h2 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_2_re) : $signed(
    _GEN_527); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_529 = 4'h3 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_3_re) : $signed(
    _GEN_528); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_530 = 4'h4 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_4_re) : $signed(
    _GEN_529); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_531 = 4'h5 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_5_re) : $signed(
    _GEN_530); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_532 = 4'h6 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_6_re) : $signed(
    _GEN_531); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_533 = 4'h7 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_7_re) : $signed(
    _GEN_532); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_534 = 4'h8 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_8_re) : $signed(
    _GEN_533); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_535 = 4'h9 == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_9_re) : $signed(
    _GEN_534); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_536 = 4'ha == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_10_re) : $signed(
    _GEN_535); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_537 = 4'hb == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_11_re) : $signed(
    _GEN_536); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_538 = 4'hc == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_12_re) : $signed(
    _GEN_537); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_539 = 4'hd == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_13_re) : $signed(
    _GEN_538); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_540 = 4'he == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_14_re) : $signed(
    _GEN_539); // @[Cholesky_V1.scala 158:{55,55}]
  wire [63:0] _GEN_541 = 4'hf == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(matrix_comp_reg_15_re) : $signed(
    _GEN_540); // @[Cholesky_V1.scala 158:{55,55}]
  wire [3:0] _GEN_544 = cholesky_comp_unit_io_valid ? 4'h3 : comp_status; // @[Cholesky_V1.scala 169:41 170:21 129:34]
  wire [31:0] _matrix_comp_reg_0_T_1 = 32'h0 - point_index; // @[Cholesky_V1.scala 177:79]
  wire [34:0] _matrix_comp_reg_0_T_2 = _matrix_comp_reg_0_T_1 * 3'h4; // @[Cholesky_V1.scala 177:93]
  wire [34:0] _GEN_1376 = {{3'd0}, _matrix_comp_reg_0_T_1}; // @[Cholesky_V1.scala 177:99]
  wire [34:0] _matrix_comp_reg_0_T_6 = _matrix_comp_reg_0_T_2 + _GEN_1376; // @[Cholesky_V1.scala 177:99]
  wire [63:0] _GEN_545 = cholesky_comp_unit_io_matrixOut_0_im; // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_546 = 4'h1 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_im) : $signed(
    _GEN_545); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_547 = 4'h2 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_im) : $signed(
    _GEN_546); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_548 = 4'h3 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_im) : $signed(
    _GEN_547); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_549 = 4'h4 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_im) : $signed(
    _GEN_548); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_550 = 4'h5 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_im) : $signed(
    _GEN_549); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_551 = 4'h6 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_im) : $signed(
    _GEN_550); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_552 = 4'h7 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_im) : $signed(
    _GEN_551); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_553 = 4'h8 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_im) : $signed(
    _GEN_552); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_554 = 4'h9 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_im) : $signed(
    _GEN_553); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_555 = 4'ha == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_im) : $signed(
    _GEN_554); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_556 = 4'hb == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_im) : $signed(
    _GEN_555); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_557 = 4'hc == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_im) : $signed(
    _GEN_556); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_558 = 4'hd == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_im) : $signed(
    _GEN_557); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_559 = 4'he == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_im) : $signed(
    _GEN_558); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_560 = 4'hf == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_im) : $signed(
    _GEN_559); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_561 = cholesky_comp_unit_io_matrixOut_0_re; // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_562 = 4'h1 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_re) : $signed(
    _GEN_561); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_563 = 4'h2 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_re) : $signed(
    _GEN_562); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_564 = 4'h3 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_re) : $signed(
    _GEN_563); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_565 = 4'h4 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_re) : $signed(
    _GEN_564); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_566 = 4'h5 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_re) : $signed(
    _GEN_565); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_567 = 4'h6 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_re) : $signed(
    _GEN_566); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_568 = 4'h7 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_re) : $signed(
    _GEN_567); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_569 = 4'h8 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_re) : $signed(
    _GEN_568); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_570 = 4'h9 == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_re) : $signed(
    _GEN_569); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_571 = 4'ha == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_re) : $signed(
    _GEN_570); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_572 = 4'hb == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_re) : $signed(
    _GEN_571); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_573 = 4'hc == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_re) : $signed(
    _GEN_572); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_574 = 4'hd == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_re) : $signed(
    _GEN_573); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_575 = 4'he == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_re) : $signed(
    _GEN_574); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_576 = 4'hf == _matrix_comp_reg_0_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_re) : $signed(
    _GEN_575); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_577 = 32'h0 >= point_index & 32'h0 >= point_index ? $signed(_GEN_560) : $signed(matrix_comp_reg_0_im)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [63:0] _GEN_578 = 32'h0 >= point_index & 32'h0 >= point_index ? $signed(_GEN_576) : $signed(matrix_comp_reg_0_re)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [31:0] _matrix_comp_reg_1_T_4 = 32'h1 - point_index; // @[Cholesky_V1.scala 177:105]
  wire [34:0] _GEN_1377 = {{3'd0}, _matrix_comp_reg_1_T_4}; // @[Cholesky_V1.scala 177:99]
  wire [34:0] _matrix_comp_reg_1_T_6 = _matrix_comp_reg_0_T_2 + _GEN_1377; // @[Cholesky_V1.scala 177:99]
  wire [63:0] _GEN_580 = 4'h1 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_im) : $signed(
    _GEN_545); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_581 = 4'h2 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_im) : $signed(
    _GEN_580); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_582 = 4'h3 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_im) : $signed(
    _GEN_581); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_583 = 4'h4 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_im) : $signed(
    _GEN_582); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_584 = 4'h5 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_im) : $signed(
    _GEN_583); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_585 = 4'h6 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_im) : $signed(
    _GEN_584); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_586 = 4'h7 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_im) : $signed(
    _GEN_585); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_587 = 4'h8 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_im) : $signed(
    _GEN_586); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_588 = 4'h9 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_im) : $signed(
    _GEN_587); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_589 = 4'ha == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_im) : $signed(
    _GEN_588); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_590 = 4'hb == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_im) : $signed(
    _GEN_589); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_591 = 4'hc == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_im) : $signed(
    _GEN_590); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_592 = 4'hd == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_im) : $signed(
    _GEN_591); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_593 = 4'he == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_im) : $signed(
    _GEN_592); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_594 = 4'hf == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_im) : $signed(
    _GEN_593); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_596 = 4'h1 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_re) : $signed(
    _GEN_561); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_597 = 4'h2 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_re) : $signed(
    _GEN_596); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_598 = 4'h3 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_re) : $signed(
    _GEN_597); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_599 = 4'h4 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_re) : $signed(
    _GEN_598); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_600 = 4'h5 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_re) : $signed(
    _GEN_599); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_601 = 4'h6 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_re) : $signed(
    _GEN_600); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_602 = 4'h7 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_re) : $signed(
    _GEN_601); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_603 = 4'h8 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_re) : $signed(
    _GEN_602); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_604 = 4'h9 == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_re) : $signed(
    _GEN_603); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_605 = 4'ha == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_re) : $signed(
    _GEN_604); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_606 = 4'hb == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_re) : $signed(
    _GEN_605); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_607 = 4'hc == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_re) : $signed(
    _GEN_606); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_608 = 4'hd == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_re) : $signed(
    _GEN_607); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_609 = 4'he == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_re) : $signed(
    _GEN_608); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_610 = 4'hf == _matrix_comp_reg_1_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_re) : $signed(
    _GEN_609); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_611 = 32'h0 >= point_index & 32'h1 >= point_index ? $signed(_GEN_594) : $signed(matrix_comp_reg_1_im)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [63:0] _GEN_612 = 32'h0 >= point_index & 32'h1 >= point_index ? $signed(_GEN_610) : $signed(matrix_comp_reg_1_re)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [31:0] _matrix_comp_reg_2_T_4 = 32'h2 - point_index; // @[Cholesky_V1.scala 177:105]
  wire [34:0] _GEN_1378 = {{3'd0}, _matrix_comp_reg_2_T_4}; // @[Cholesky_V1.scala 177:99]
  wire [34:0] _matrix_comp_reg_2_T_6 = _matrix_comp_reg_0_T_2 + _GEN_1378; // @[Cholesky_V1.scala 177:99]
  wire [63:0] _GEN_614 = 4'h1 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_im) : $signed(
    _GEN_545); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_615 = 4'h2 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_im) : $signed(
    _GEN_614); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_616 = 4'h3 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_im) : $signed(
    _GEN_615); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_617 = 4'h4 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_im) : $signed(
    _GEN_616); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_618 = 4'h5 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_im) : $signed(
    _GEN_617); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_619 = 4'h6 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_im) : $signed(
    _GEN_618); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_620 = 4'h7 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_im) : $signed(
    _GEN_619); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_621 = 4'h8 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_im) : $signed(
    _GEN_620); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_622 = 4'h9 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_im) : $signed(
    _GEN_621); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_623 = 4'ha == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_im) : $signed(
    _GEN_622); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_624 = 4'hb == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_im) : $signed(
    _GEN_623); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_625 = 4'hc == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_im) : $signed(
    _GEN_624); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_626 = 4'hd == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_im) : $signed(
    _GEN_625); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_627 = 4'he == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_im) : $signed(
    _GEN_626); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_628 = 4'hf == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_im) : $signed(
    _GEN_627); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_630 = 4'h1 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_re) : $signed(
    _GEN_561); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_631 = 4'h2 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_re) : $signed(
    _GEN_630); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_632 = 4'h3 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_re) : $signed(
    _GEN_631); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_633 = 4'h4 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_re) : $signed(
    _GEN_632); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_634 = 4'h5 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_re) : $signed(
    _GEN_633); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_635 = 4'h6 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_re) : $signed(
    _GEN_634); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_636 = 4'h7 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_re) : $signed(
    _GEN_635); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_637 = 4'h8 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_re) : $signed(
    _GEN_636); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_638 = 4'h9 == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_re) : $signed(
    _GEN_637); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_639 = 4'ha == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_re) : $signed(
    _GEN_638); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_640 = 4'hb == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_re) : $signed(
    _GEN_639); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_641 = 4'hc == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_re) : $signed(
    _GEN_640); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_642 = 4'hd == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_re) : $signed(
    _GEN_641); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_643 = 4'he == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_re) : $signed(
    _GEN_642); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_644 = 4'hf == _matrix_comp_reg_2_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_re) : $signed(
    _GEN_643); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_645 = 32'h0 >= point_index & 32'h2 >= point_index ? $signed(_GEN_628) : $signed(matrix_comp_reg_2_im)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [63:0] _GEN_646 = 32'h0 >= point_index & 32'h2 >= point_index ? $signed(_GEN_644) : $signed(matrix_comp_reg_2_re)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [31:0] _matrix_comp_reg_3_T_4 = 32'h3 - point_index; // @[Cholesky_V1.scala 177:105]
  wire [34:0] _GEN_1379 = {{3'd0}, _matrix_comp_reg_3_T_4}; // @[Cholesky_V1.scala 177:99]
  wire [34:0] _matrix_comp_reg_3_T_6 = _matrix_comp_reg_0_T_2 + _GEN_1379; // @[Cholesky_V1.scala 177:99]
  wire [63:0] _GEN_648 = 4'h1 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_im) : $signed(
    _GEN_545); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_649 = 4'h2 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_im) : $signed(
    _GEN_648); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_650 = 4'h3 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_im) : $signed(
    _GEN_649); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_651 = 4'h4 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_im) : $signed(
    _GEN_650); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_652 = 4'h5 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_im) : $signed(
    _GEN_651); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_653 = 4'h6 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_im) : $signed(
    _GEN_652); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_654 = 4'h7 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_im) : $signed(
    _GEN_653); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_655 = 4'h8 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_im) : $signed(
    _GEN_654); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_656 = 4'h9 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_im) : $signed(
    _GEN_655); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_657 = 4'ha == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_im) : $signed(
    _GEN_656); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_658 = 4'hb == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_im) : $signed(
    _GEN_657); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_659 = 4'hc == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_im) : $signed(
    _GEN_658); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_660 = 4'hd == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_im) : $signed(
    _GEN_659); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_661 = 4'he == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_im) : $signed(
    _GEN_660); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_662 = 4'hf == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_im) : $signed(
    _GEN_661); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_664 = 4'h1 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_re) : $signed(
    _GEN_561); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_665 = 4'h2 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_re) : $signed(
    _GEN_664); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_666 = 4'h3 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_re) : $signed(
    _GEN_665); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_667 = 4'h4 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_re) : $signed(
    _GEN_666); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_668 = 4'h5 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_re) : $signed(
    _GEN_667); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_669 = 4'h6 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_re) : $signed(
    _GEN_668); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_670 = 4'h7 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_re) : $signed(
    _GEN_669); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_671 = 4'h8 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_re) : $signed(
    _GEN_670); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_672 = 4'h9 == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_re) : $signed(
    _GEN_671); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_673 = 4'ha == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_re) : $signed(
    _GEN_672); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_674 = 4'hb == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_re) : $signed(
    _GEN_673); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_675 = 4'hc == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_re) : $signed(
    _GEN_674); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_676 = 4'hd == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_re) : $signed(
    _GEN_675); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_677 = 4'he == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_re) : $signed(
    _GEN_676); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_678 = 4'hf == _matrix_comp_reg_3_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_re) : $signed(
    _GEN_677); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_679 = 32'h0 >= point_index & 32'h3 >= point_index ? $signed(_GEN_662) : $signed(matrix_comp_reg_3_im)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [63:0] _GEN_680 = 32'h0 >= point_index & 32'h3 >= point_index ? $signed(_GEN_678) : $signed(matrix_comp_reg_3_re)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [34:0] _matrix_comp_reg_4_T_2 = _matrix_comp_reg_1_T_4 * 3'h4; // @[Cholesky_V1.scala 177:93]
  wire [34:0] _matrix_comp_reg_4_T_6 = _matrix_comp_reg_4_T_2 + _GEN_1376; // @[Cholesky_V1.scala 177:99]
  wire [63:0] _GEN_682 = 4'h1 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_im) : $signed(
    _GEN_545); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_683 = 4'h2 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_im) : $signed(
    _GEN_682); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_684 = 4'h3 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_im) : $signed(
    _GEN_683); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_685 = 4'h4 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_im) : $signed(
    _GEN_684); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_686 = 4'h5 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_im) : $signed(
    _GEN_685); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_687 = 4'h6 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_im) : $signed(
    _GEN_686); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_688 = 4'h7 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_im) : $signed(
    _GEN_687); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_689 = 4'h8 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_im) : $signed(
    _GEN_688); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_690 = 4'h9 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_im) : $signed(
    _GEN_689); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_691 = 4'ha == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_im) : $signed(
    _GEN_690); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_692 = 4'hb == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_im) : $signed(
    _GEN_691); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_693 = 4'hc == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_im) : $signed(
    _GEN_692); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_694 = 4'hd == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_im) : $signed(
    _GEN_693); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_695 = 4'he == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_im) : $signed(
    _GEN_694); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_696 = 4'hf == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_im) : $signed(
    _GEN_695); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_698 = 4'h1 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_re) : $signed(
    _GEN_561); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_699 = 4'h2 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_re) : $signed(
    _GEN_698); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_700 = 4'h3 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_re) : $signed(
    _GEN_699); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_701 = 4'h4 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_re) : $signed(
    _GEN_700); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_702 = 4'h5 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_re) : $signed(
    _GEN_701); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_703 = 4'h6 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_re) : $signed(
    _GEN_702); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_704 = 4'h7 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_re) : $signed(
    _GEN_703); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_705 = 4'h8 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_re) : $signed(
    _GEN_704); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_706 = 4'h9 == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_re) : $signed(
    _GEN_705); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_707 = 4'ha == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_re) : $signed(
    _GEN_706); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_708 = 4'hb == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_re) : $signed(
    _GEN_707); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_709 = 4'hc == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_re) : $signed(
    _GEN_708); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_710 = 4'hd == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_re) : $signed(
    _GEN_709); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_711 = 4'he == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_re) : $signed(
    _GEN_710); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_712 = 4'hf == _matrix_comp_reg_4_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_re) : $signed(
    _GEN_711); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_713 = 32'h1 >= point_index & 32'h0 >= point_index ? $signed(_GEN_696) : $signed(matrix_comp_reg_4_im)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [63:0] _GEN_714 = 32'h1 >= point_index & 32'h0 >= point_index ? $signed(_GEN_712) : $signed(matrix_comp_reg_4_re)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [34:0] _matrix_comp_reg_5_T_6 = _matrix_comp_reg_4_T_2 + _GEN_1377; // @[Cholesky_V1.scala 177:99]
  wire [63:0] _GEN_716 = 4'h1 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_im) : $signed(
    _GEN_545); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_717 = 4'h2 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_im) : $signed(
    _GEN_716); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_718 = 4'h3 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_im) : $signed(
    _GEN_717); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_719 = 4'h4 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_im) : $signed(
    _GEN_718); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_720 = 4'h5 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_im) : $signed(
    _GEN_719); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_721 = 4'h6 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_im) : $signed(
    _GEN_720); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_722 = 4'h7 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_im) : $signed(
    _GEN_721); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_723 = 4'h8 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_im) : $signed(
    _GEN_722); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_724 = 4'h9 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_im) : $signed(
    _GEN_723); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_725 = 4'ha == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_im) : $signed(
    _GEN_724); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_726 = 4'hb == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_im) : $signed(
    _GEN_725); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_727 = 4'hc == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_im) : $signed(
    _GEN_726); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_728 = 4'hd == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_im) : $signed(
    _GEN_727); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_729 = 4'he == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_im) : $signed(
    _GEN_728); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_730 = 4'hf == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_im) : $signed(
    _GEN_729); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_732 = 4'h1 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_re) : $signed(
    _GEN_561); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_733 = 4'h2 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_re) : $signed(
    _GEN_732); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_734 = 4'h3 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_re) : $signed(
    _GEN_733); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_735 = 4'h4 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_re) : $signed(
    _GEN_734); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_736 = 4'h5 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_re) : $signed(
    _GEN_735); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_737 = 4'h6 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_re) : $signed(
    _GEN_736); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_738 = 4'h7 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_re) : $signed(
    _GEN_737); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_739 = 4'h8 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_re) : $signed(
    _GEN_738); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_740 = 4'h9 == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_re) : $signed(
    _GEN_739); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_741 = 4'ha == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_re) : $signed(
    _GEN_740); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_742 = 4'hb == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_re) : $signed(
    _GEN_741); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_743 = 4'hc == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_re) : $signed(
    _GEN_742); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_744 = 4'hd == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_re) : $signed(
    _GEN_743); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_745 = 4'he == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_re) : $signed(
    _GEN_744); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_746 = 4'hf == _matrix_comp_reg_5_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_re) : $signed(
    _GEN_745); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_747 = 32'h1 >= point_index & 32'h1 >= point_index ? $signed(_GEN_730) : $signed(matrix_comp_reg_5_im)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [63:0] _GEN_748 = 32'h1 >= point_index & 32'h1 >= point_index ? $signed(_GEN_746) : $signed(matrix_comp_reg_5_re)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [34:0] _matrix_comp_reg_6_T_6 = _matrix_comp_reg_4_T_2 + _GEN_1378; // @[Cholesky_V1.scala 177:99]
  wire [63:0] _GEN_750 = 4'h1 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_im) : $signed(
    _GEN_545); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_751 = 4'h2 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_im) : $signed(
    _GEN_750); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_752 = 4'h3 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_im) : $signed(
    _GEN_751); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_753 = 4'h4 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_im) : $signed(
    _GEN_752); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_754 = 4'h5 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_im) : $signed(
    _GEN_753); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_755 = 4'h6 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_im) : $signed(
    _GEN_754); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_756 = 4'h7 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_im) : $signed(
    _GEN_755); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_757 = 4'h8 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_im) : $signed(
    _GEN_756); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_758 = 4'h9 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_im) : $signed(
    _GEN_757); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_759 = 4'ha == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_im) : $signed(
    _GEN_758); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_760 = 4'hb == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_im) : $signed(
    _GEN_759); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_761 = 4'hc == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_im) : $signed(
    _GEN_760); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_762 = 4'hd == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_im) : $signed(
    _GEN_761); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_763 = 4'he == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_im) : $signed(
    _GEN_762); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_764 = 4'hf == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_im) : $signed(
    _GEN_763); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_766 = 4'h1 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_re) : $signed(
    _GEN_561); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_767 = 4'h2 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_re) : $signed(
    _GEN_766); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_768 = 4'h3 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_re) : $signed(
    _GEN_767); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_769 = 4'h4 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_re) : $signed(
    _GEN_768); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_770 = 4'h5 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_re) : $signed(
    _GEN_769); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_771 = 4'h6 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_re) : $signed(
    _GEN_770); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_772 = 4'h7 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_re) : $signed(
    _GEN_771); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_773 = 4'h8 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_re) : $signed(
    _GEN_772); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_774 = 4'h9 == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_re) : $signed(
    _GEN_773); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_775 = 4'ha == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_re) : $signed(
    _GEN_774); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_776 = 4'hb == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_re) : $signed(
    _GEN_775); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_777 = 4'hc == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_re) : $signed(
    _GEN_776); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_778 = 4'hd == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_re) : $signed(
    _GEN_777); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_779 = 4'he == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_re) : $signed(
    _GEN_778); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_780 = 4'hf == _matrix_comp_reg_6_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_re) : $signed(
    _GEN_779); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_781 = 32'h1 >= point_index & 32'h2 >= point_index ? $signed(_GEN_764) : $signed(matrix_comp_reg_6_im)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [63:0] _GEN_782 = 32'h1 >= point_index & 32'h2 >= point_index ? $signed(_GEN_780) : $signed(matrix_comp_reg_6_re)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [34:0] _matrix_comp_reg_7_T_6 = _matrix_comp_reg_4_T_2 + _GEN_1379; // @[Cholesky_V1.scala 177:99]
  wire [63:0] _GEN_784 = 4'h1 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_im) : $signed(
    _GEN_545); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_785 = 4'h2 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_im) : $signed(
    _GEN_784); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_786 = 4'h3 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_im) : $signed(
    _GEN_785); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_787 = 4'h4 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_im) : $signed(
    _GEN_786); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_788 = 4'h5 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_im) : $signed(
    _GEN_787); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_789 = 4'h6 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_im) : $signed(
    _GEN_788); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_790 = 4'h7 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_im) : $signed(
    _GEN_789); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_791 = 4'h8 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_im) : $signed(
    _GEN_790); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_792 = 4'h9 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_im) : $signed(
    _GEN_791); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_793 = 4'ha == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_im) : $signed(
    _GEN_792); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_794 = 4'hb == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_im) : $signed(
    _GEN_793); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_795 = 4'hc == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_im) : $signed(
    _GEN_794); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_796 = 4'hd == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_im) : $signed(
    _GEN_795); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_797 = 4'he == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_im) : $signed(
    _GEN_796); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_798 = 4'hf == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_im) : $signed(
    _GEN_797); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_800 = 4'h1 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_re) : $signed(
    _GEN_561); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_801 = 4'h2 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_re) : $signed(
    _GEN_800); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_802 = 4'h3 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_re) : $signed(
    _GEN_801); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_803 = 4'h4 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_re) : $signed(
    _GEN_802); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_804 = 4'h5 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_re) : $signed(
    _GEN_803); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_805 = 4'h6 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_re) : $signed(
    _GEN_804); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_806 = 4'h7 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_re) : $signed(
    _GEN_805); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_807 = 4'h8 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_re) : $signed(
    _GEN_806); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_808 = 4'h9 == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_re) : $signed(
    _GEN_807); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_809 = 4'ha == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_re) : $signed(
    _GEN_808); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_810 = 4'hb == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_re) : $signed(
    _GEN_809); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_811 = 4'hc == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_re) : $signed(
    _GEN_810); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_812 = 4'hd == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_re) : $signed(
    _GEN_811); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_813 = 4'he == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_re) : $signed(
    _GEN_812); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_814 = 4'hf == _matrix_comp_reg_7_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_re) : $signed(
    _GEN_813); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_815 = 32'h1 >= point_index & 32'h3 >= point_index ? $signed(_GEN_798) : $signed(matrix_comp_reg_7_im)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [63:0] _GEN_816 = 32'h1 >= point_index & 32'h3 >= point_index ? $signed(_GEN_814) : $signed(matrix_comp_reg_7_re)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [34:0] _matrix_comp_reg_8_T_2 = _matrix_comp_reg_2_T_4 * 3'h4; // @[Cholesky_V1.scala 177:93]
  wire [34:0] _matrix_comp_reg_8_T_6 = _matrix_comp_reg_8_T_2 + _GEN_1376; // @[Cholesky_V1.scala 177:99]
  wire [63:0] _GEN_818 = 4'h1 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_im) : $signed(
    _GEN_545); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_819 = 4'h2 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_im) : $signed(
    _GEN_818); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_820 = 4'h3 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_im) : $signed(
    _GEN_819); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_821 = 4'h4 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_im) : $signed(
    _GEN_820); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_822 = 4'h5 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_im) : $signed(
    _GEN_821); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_823 = 4'h6 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_im) : $signed(
    _GEN_822); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_824 = 4'h7 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_im) : $signed(
    _GEN_823); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_825 = 4'h8 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_im) : $signed(
    _GEN_824); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_826 = 4'h9 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_im) : $signed(
    _GEN_825); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_827 = 4'ha == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_im) : $signed(
    _GEN_826); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_828 = 4'hb == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_im) : $signed(
    _GEN_827); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_829 = 4'hc == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_im) : $signed(
    _GEN_828); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_830 = 4'hd == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_im) : $signed(
    _GEN_829); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_831 = 4'he == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_im) : $signed(
    _GEN_830); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_832 = 4'hf == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_im) : $signed(
    _GEN_831); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_834 = 4'h1 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_re) : $signed(
    _GEN_561); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_835 = 4'h2 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_re) : $signed(
    _GEN_834); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_836 = 4'h3 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_re) : $signed(
    _GEN_835); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_837 = 4'h4 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_re) : $signed(
    _GEN_836); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_838 = 4'h5 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_re) : $signed(
    _GEN_837); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_839 = 4'h6 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_re) : $signed(
    _GEN_838); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_840 = 4'h7 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_re) : $signed(
    _GEN_839); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_841 = 4'h8 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_re) : $signed(
    _GEN_840); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_842 = 4'h9 == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_re) : $signed(
    _GEN_841); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_843 = 4'ha == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_re) : $signed(
    _GEN_842); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_844 = 4'hb == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_re) : $signed(
    _GEN_843); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_845 = 4'hc == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_re) : $signed(
    _GEN_844); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_846 = 4'hd == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_re) : $signed(
    _GEN_845); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_847 = 4'he == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_re) : $signed(
    _GEN_846); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_848 = 4'hf == _matrix_comp_reg_8_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_re) : $signed(
    _GEN_847); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_849 = 32'h2 >= point_index & 32'h0 >= point_index ? $signed(_GEN_832) : $signed(matrix_comp_reg_8_im)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [63:0] _GEN_850 = 32'h2 >= point_index & 32'h0 >= point_index ? $signed(_GEN_848) : $signed(matrix_comp_reg_8_re)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [34:0] _matrix_comp_reg_9_T_6 = _matrix_comp_reg_8_T_2 + _GEN_1377; // @[Cholesky_V1.scala 177:99]
  wire [63:0] _GEN_852 = 4'h1 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_im) : $signed(
    _GEN_545); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_853 = 4'h2 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_im) : $signed(
    _GEN_852); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_854 = 4'h3 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_im) : $signed(
    _GEN_853); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_855 = 4'h4 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_im) : $signed(
    _GEN_854); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_856 = 4'h5 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_im) : $signed(
    _GEN_855); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_857 = 4'h6 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_im) : $signed(
    _GEN_856); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_858 = 4'h7 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_im) : $signed(
    _GEN_857); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_859 = 4'h8 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_im) : $signed(
    _GEN_858); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_860 = 4'h9 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_im) : $signed(
    _GEN_859); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_861 = 4'ha == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_im) : $signed(
    _GEN_860); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_862 = 4'hb == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_im) : $signed(
    _GEN_861); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_863 = 4'hc == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_im) : $signed(
    _GEN_862); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_864 = 4'hd == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_im) : $signed(
    _GEN_863); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_865 = 4'he == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_im) : $signed(
    _GEN_864); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_866 = 4'hf == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_im) : $signed(
    _GEN_865); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_868 = 4'h1 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_re) : $signed(
    _GEN_561); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_869 = 4'h2 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_re) : $signed(
    _GEN_868); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_870 = 4'h3 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_re) : $signed(
    _GEN_869); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_871 = 4'h4 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_re) : $signed(
    _GEN_870); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_872 = 4'h5 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_re) : $signed(
    _GEN_871); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_873 = 4'h6 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_re) : $signed(
    _GEN_872); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_874 = 4'h7 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_re) : $signed(
    _GEN_873); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_875 = 4'h8 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_re) : $signed(
    _GEN_874); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_876 = 4'h9 == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_re) : $signed(
    _GEN_875); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_877 = 4'ha == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_re) : $signed(
    _GEN_876); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_878 = 4'hb == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_re) : $signed(
    _GEN_877); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_879 = 4'hc == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_re) : $signed(
    _GEN_878); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_880 = 4'hd == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_re) : $signed(
    _GEN_879); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_881 = 4'he == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_re) : $signed(
    _GEN_880); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_882 = 4'hf == _matrix_comp_reg_9_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_re) : $signed(
    _GEN_881); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_883 = 32'h2 >= point_index & 32'h1 >= point_index ? $signed(_GEN_866) : $signed(matrix_comp_reg_9_im)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [63:0] _GEN_884 = 32'h2 >= point_index & 32'h1 >= point_index ? $signed(_GEN_882) : $signed(matrix_comp_reg_9_re)
    ; // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [34:0] _matrix_comp_reg_10_T_6 = _matrix_comp_reg_8_T_2 + _GEN_1378; // @[Cholesky_V1.scala 177:99]
  wire [63:0] _GEN_886 = 4'h1 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_im) : $signed(
    _GEN_545); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_887 = 4'h2 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_im) : $signed(
    _GEN_886); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_888 = 4'h3 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_im) : $signed(
    _GEN_887); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_889 = 4'h4 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_im) : $signed(
    _GEN_888); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_890 = 4'h5 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_im) : $signed(
    _GEN_889); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_891 = 4'h6 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_im) : $signed(
    _GEN_890); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_892 = 4'h7 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_im) : $signed(
    _GEN_891); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_893 = 4'h8 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_im) : $signed(
    _GEN_892); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_894 = 4'h9 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_im) : $signed(
    _GEN_893); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_895 = 4'ha == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_im) :
    $signed(_GEN_894); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_896 = 4'hb == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_im) :
    $signed(_GEN_895); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_897 = 4'hc == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_im) :
    $signed(_GEN_896); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_898 = 4'hd == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_im) :
    $signed(_GEN_897); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_899 = 4'he == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_im) :
    $signed(_GEN_898); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_900 = 4'hf == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_im) :
    $signed(_GEN_899); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_902 = 4'h1 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_re) : $signed(
    _GEN_561); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_903 = 4'h2 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_re) : $signed(
    _GEN_902); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_904 = 4'h3 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_re) : $signed(
    _GEN_903); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_905 = 4'h4 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_re) : $signed(
    _GEN_904); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_906 = 4'h5 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_re) : $signed(
    _GEN_905); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_907 = 4'h6 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_re) : $signed(
    _GEN_906); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_908 = 4'h7 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_re) : $signed(
    _GEN_907); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_909 = 4'h8 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_re) : $signed(
    _GEN_908); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_910 = 4'h9 == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_re) : $signed(
    _GEN_909); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_911 = 4'ha == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_re) :
    $signed(_GEN_910); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_912 = 4'hb == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_re) :
    $signed(_GEN_911); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_913 = 4'hc == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_re) :
    $signed(_GEN_912); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_914 = 4'hd == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_re) :
    $signed(_GEN_913); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_915 = 4'he == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_re) :
    $signed(_GEN_914); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_916 = 4'hf == _matrix_comp_reg_10_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_re) :
    $signed(_GEN_915); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_917 = 32'h2 >= point_index & 32'h2 >= point_index ? $signed(_GEN_900) : $signed(matrix_comp_reg_10_im
    ); // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [63:0] _GEN_918 = 32'h2 >= point_index & 32'h2 >= point_index ? $signed(_GEN_916) : $signed(matrix_comp_reg_10_re
    ); // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [34:0] _matrix_comp_reg_11_T_6 = _matrix_comp_reg_8_T_2 + _GEN_1379; // @[Cholesky_V1.scala 177:99]
  wire [63:0] _GEN_920 = 4'h1 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_im) : $signed(
    _GEN_545); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_921 = 4'h2 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_im) : $signed(
    _GEN_920); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_922 = 4'h3 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_im) : $signed(
    _GEN_921); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_923 = 4'h4 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_im) : $signed(
    _GEN_922); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_924 = 4'h5 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_im) : $signed(
    _GEN_923); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_925 = 4'h6 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_im) : $signed(
    _GEN_924); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_926 = 4'h7 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_im) : $signed(
    _GEN_925); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_927 = 4'h8 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_im) : $signed(
    _GEN_926); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_928 = 4'h9 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_im) : $signed(
    _GEN_927); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_929 = 4'ha == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_im) :
    $signed(_GEN_928); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_930 = 4'hb == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_im) :
    $signed(_GEN_929); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_931 = 4'hc == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_im) :
    $signed(_GEN_930); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_932 = 4'hd == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_im) :
    $signed(_GEN_931); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_933 = 4'he == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_im) :
    $signed(_GEN_932); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_934 = 4'hf == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_im) :
    $signed(_GEN_933); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_936 = 4'h1 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_re) : $signed(
    _GEN_561); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_937 = 4'h2 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_re) : $signed(
    _GEN_936); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_938 = 4'h3 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_re) : $signed(
    _GEN_937); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_939 = 4'h4 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_re) : $signed(
    _GEN_938); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_940 = 4'h5 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_re) : $signed(
    _GEN_939); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_941 = 4'h6 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_re) : $signed(
    _GEN_940); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_942 = 4'h7 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_re) : $signed(
    _GEN_941); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_943 = 4'h8 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_re) : $signed(
    _GEN_942); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_944 = 4'h9 == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_re) : $signed(
    _GEN_943); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_945 = 4'ha == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_re) :
    $signed(_GEN_944); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_946 = 4'hb == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_re) :
    $signed(_GEN_945); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_947 = 4'hc == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_re) :
    $signed(_GEN_946); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_948 = 4'hd == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_re) :
    $signed(_GEN_947); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_949 = 4'he == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_re) :
    $signed(_GEN_948); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_950 = 4'hf == _matrix_comp_reg_11_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_re) :
    $signed(_GEN_949); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_951 = 32'h2 >= point_index & 32'h3 >= point_index ? $signed(_GEN_934) : $signed(matrix_comp_reg_11_im
    ); // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [63:0] _GEN_952 = 32'h2 >= point_index & 32'h3 >= point_index ? $signed(_GEN_950) : $signed(matrix_comp_reg_11_re
    ); // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [34:0] _matrix_comp_reg_12_T_2 = _matrix_comp_reg_3_T_4 * 3'h4; // @[Cholesky_V1.scala 177:93]
  wire [34:0] _matrix_comp_reg_12_T_6 = _matrix_comp_reg_12_T_2 + _GEN_1376; // @[Cholesky_V1.scala 177:99]
  wire [63:0] _GEN_954 = 4'h1 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_im) : $signed(
    _GEN_545); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_955 = 4'h2 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_im) : $signed(
    _GEN_954); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_956 = 4'h3 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_im) : $signed(
    _GEN_955); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_957 = 4'h4 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_im) : $signed(
    _GEN_956); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_958 = 4'h5 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_im) : $signed(
    _GEN_957); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_959 = 4'h6 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_im) : $signed(
    _GEN_958); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_960 = 4'h7 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_im) : $signed(
    _GEN_959); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_961 = 4'h8 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_im) : $signed(
    _GEN_960); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_962 = 4'h9 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_im) : $signed(
    _GEN_961); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_963 = 4'ha == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_im) :
    $signed(_GEN_962); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_964 = 4'hb == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_im) :
    $signed(_GEN_963); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_965 = 4'hc == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_im) :
    $signed(_GEN_964); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_966 = 4'hd == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_im) :
    $signed(_GEN_965); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_967 = 4'he == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_im) :
    $signed(_GEN_966); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_968 = 4'hf == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_im) :
    $signed(_GEN_967); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_970 = 4'h1 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_re) : $signed(
    _GEN_561); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_971 = 4'h2 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_re) : $signed(
    _GEN_970); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_972 = 4'h3 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_re) : $signed(
    _GEN_971); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_973 = 4'h4 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_re) : $signed(
    _GEN_972); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_974 = 4'h5 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_re) : $signed(
    _GEN_973); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_975 = 4'h6 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_re) : $signed(
    _GEN_974); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_976 = 4'h7 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_re) : $signed(
    _GEN_975); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_977 = 4'h8 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_re) : $signed(
    _GEN_976); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_978 = 4'h9 == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_re) : $signed(
    _GEN_977); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_979 = 4'ha == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_re) :
    $signed(_GEN_978); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_980 = 4'hb == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_re) :
    $signed(_GEN_979); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_981 = 4'hc == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_re) :
    $signed(_GEN_980); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_982 = 4'hd == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_re) :
    $signed(_GEN_981); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_983 = 4'he == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_re) :
    $signed(_GEN_982); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_984 = 4'hf == _matrix_comp_reg_12_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_re) :
    $signed(_GEN_983); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_985 = 32'h3 >= point_index & 32'h0 >= point_index ? $signed(_GEN_968) : $signed(matrix_comp_reg_12_im
    ); // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [63:0] _GEN_986 = 32'h3 >= point_index & 32'h0 >= point_index ? $signed(_GEN_984) : $signed(matrix_comp_reg_12_re
    ); // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [34:0] _matrix_comp_reg_13_T_6 = _matrix_comp_reg_12_T_2 + _GEN_1377; // @[Cholesky_V1.scala 177:99]
  wire [63:0] _GEN_988 = 4'h1 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_im) : $signed(
    _GEN_545); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_989 = 4'h2 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_im) : $signed(
    _GEN_988); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_990 = 4'h3 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_im) : $signed(
    _GEN_989); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_991 = 4'h4 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_im) : $signed(
    _GEN_990); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_992 = 4'h5 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_im) : $signed(
    _GEN_991); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_993 = 4'h6 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_im) : $signed(
    _GEN_992); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_994 = 4'h7 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_im) : $signed(
    _GEN_993); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_995 = 4'h8 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_im) : $signed(
    _GEN_994); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_996 = 4'h9 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_im) : $signed(
    _GEN_995); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_997 = 4'ha == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_im) :
    $signed(_GEN_996); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_998 = 4'hb == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_im) :
    $signed(_GEN_997); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_999 = 4'hc == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_im) :
    $signed(_GEN_998); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1000 = 4'hd == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_im) :
    $signed(_GEN_999); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1001 = 4'he == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_im) :
    $signed(_GEN_1000); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1002 = 4'hf == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_im) :
    $signed(_GEN_1001); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1004 = 4'h1 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_re) :
    $signed(_GEN_561); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1005 = 4'h2 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_re) :
    $signed(_GEN_1004); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1006 = 4'h3 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_re) :
    $signed(_GEN_1005); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1007 = 4'h4 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_re) :
    $signed(_GEN_1006); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1008 = 4'h5 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_re) :
    $signed(_GEN_1007); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1009 = 4'h6 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_re) :
    $signed(_GEN_1008); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1010 = 4'h7 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_re) :
    $signed(_GEN_1009); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1011 = 4'h8 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_re) :
    $signed(_GEN_1010); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1012 = 4'h9 == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_re) :
    $signed(_GEN_1011); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1013 = 4'ha == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_re) :
    $signed(_GEN_1012); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1014 = 4'hb == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_re) :
    $signed(_GEN_1013); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1015 = 4'hc == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_re) :
    $signed(_GEN_1014); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1016 = 4'hd == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_re) :
    $signed(_GEN_1015); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1017 = 4'he == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_re) :
    $signed(_GEN_1016); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1018 = 4'hf == _matrix_comp_reg_13_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_re) :
    $signed(_GEN_1017); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1019 = 32'h3 >= point_index & 32'h1 >= point_index ? $signed(_GEN_1002) : $signed(
    matrix_comp_reg_13_im); // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [63:0] _GEN_1020 = 32'h3 >= point_index & 32'h1 >= point_index ? $signed(_GEN_1018) : $signed(
    matrix_comp_reg_13_re); // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [34:0] _matrix_comp_reg_14_T_6 = _matrix_comp_reg_12_T_2 + _GEN_1378; // @[Cholesky_V1.scala 177:99]
  wire [63:0] _GEN_1022 = 4'h1 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_im) :
    $signed(_GEN_545); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1023 = 4'h2 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_im) :
    $signed(_GEN_1022); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1024 = 4'h3 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_im) :
    $signed(_GEN_1023); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1025 = 4'h4 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_im) :
    $signed(_GEN_1024); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1026 = 4'h5 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_im) :
    $signed(_GEN_1025); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1027 = 4'h6 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_im) :
    $signed(_GEN_1026); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1028 = 4'h7 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_im) :
    $signed(_GEN_1027); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1029 = 4'h8 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_im) :
    $signed(_GEN_1028); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1030 = 4'h9 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_im) :
    $signed(_GEN_1029); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1031 = 4'ha == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_im) :
    $signed(_GEN_1030); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1032 = 4'hb == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_im) :
    $signed(_GEN_1031); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1033 = 4'hc == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_im) :
    $signed(_GEN_1032); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1034 = 4'hd == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_im) :
    $signed(_GEN_1033); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1035 = 4'he == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_im) :
    $signed(_GEN_1034); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1036 = 4'hf == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_im) :
    $signed(_GEN_1035); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1038 = 4'h1 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_re) :
    $signed(_GEN_561); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1039 = 4'h2 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_re) :
    $signed(_GEN_1038); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1040 = 4'h3 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_re) :
    $signed(_GEN_1039); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1041 = 4'h4 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_re) :
    $signed(_GEN_1040); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1042 = 4'h5 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_re) :
    $signed(_GEN_1041); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1043 = 4'h6 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_re) :
    $signed(_GEN_1042); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1044 = 4'h7 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_re) :
    $signed(_GEN_1043); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1045 = 4'h8 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_re) :
    $signed(_GEN_1044); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1046 = 4'h9 == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_re) :
    $signed(_GEN_1045); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1047 = 4'ha == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_re) :
    $signed(_GEN_1046); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1048 = 4'hb == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_re) :
    $signed(_GEN_1047); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1049 = 4'hc == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_re) :
    $signed(_GEN_1048); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1050 = 4'hd == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_re) :
    $signed(_GEN_1049); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1051 = 4'he == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_re) :
    $signed(_GEN_1050); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1052 = 4'hf == _matrix_comp_reg_14_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_re) :
    $signed(_GEN_1051); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1053 = 32'h3 >= point_index & 32'h2 >= point_index ? $signed(_GEN_1036) : $signed(
    matrix_comp_reg_14_im); // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [63:0] _GEN_1054 = 32'h3 >= point_index & 32'h2 >= point_index ? $signed(_GEN_1052) : $signed(
    matrix_comp_reg_14_re); // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [34:0] _matrix_comp_reg_15_T_6 = _matrix_comp_reg_12_T_2 + _GEN_1379; // @[Cholesky_V1.scala 177:99]
  wire [63:0] _GEN_1056 = 4'h1 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_im) :
    $signed(_GEN_545); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1057 = 4'h2 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_im) :
    $signed(_GEN_1056); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1058 = 4'h3 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_im) :
    $signed(_GEN_1057); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1059 = 4'h4 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_im) :
    $signed(_GEN_1058); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1060 = 4'h5 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_im) :
    $signed(_GEN_1059); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1061 = 4'h6 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_im) :
    $signed(_GEN_1060); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1062 = 4'h7 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_im) :
    $signed(_GEN_1061); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1063 = 4'h8 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_im) :
    $signed(_GEN_1062); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1064 = 4'h9 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_im) :
    $signed(_GEN_1063); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1065 = 4'ha == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_im) :
    $signed(_GEN_1064); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1066 = 4'hb == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_im) :
    $signed(_GEN_1065); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1067 = 4'hc == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_im) :
    $signed(_GEN_1066); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1068 = 4'hd == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_im) :
    $signed(_GEN_1067); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1069 = 4'he == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_im) :
    $signed(_GEN_1068); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1070 = 4'hf == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_im) :
    $signed(_GEN_1069); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1072 = 4'h1 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_1_re) :
    $signed(_GEN_561); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1073 = 4'h2 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_2_re) :
    $signed(_GEN_1072); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1074 = 4'h3 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_3_re) :
    $signed(_GEN_1073); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1075 = 4'h4 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_4_re) :
    $signed(_GEN_1074); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1076 = 4'h5 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_5_re) :
    $signed(_GEN_1075); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1077 = 4'h6 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_6_re) :
    $signed(_GEN_1076); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1078 = 4'h7 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_7_re) :
    $signed(_GEN_1077); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1079 = 4'h8 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_8_re) :
    $signed(_GEN_1078); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1080 = 4'h9 == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_9_re) :
    $signed(_GEN_1079); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1081 = 4'ha == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_10_re) :
    $signed(_GEN_1080); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1082 = 4'hb == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_11_re) :
    $signed(_GEN_1081); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1083 = 4'hc == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_12_re) :
    $signed(_GEN_1082); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1084 = 4'hd == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_13_re) :
    $signed(_GEN_1083); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1085 = 4'he == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_14_re) :
    $signed(_GEN_1084); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1086 = 4'hf == _matrix_comp_reg_15_T_6[3:0] ? $signed(cholesky_comp_unit_io_matrixOut_15_re) :
    $signed(_GEN_1085); // @[Cholesky_V1.scala 177:{40,40}]
  wire [63:0] _GEN_1087 = 32'h3 >= point_index & 32'h3 >= point_index ? $signed(_GEN_1070) : $signed(
    matrix_comp_reg_15_im); // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [63:0] _GEN_1088 = 32'h3 >= point_index & 32'h3 >= point_index ? $signed(_GEN_1086) : $signed(
    matrix_comp_reg_15_re); // @[Cholesky_V1.scala 176:58 177:40 127:42]
  wire [31:0] _point_index_T_1 = point_index + 32'h1; // @[Cholesky_V1.scala 181:34]
  wire [63:0] _GEN_1089 = comp_status == 4'h3 ? $signed(_GEN_577) : $signed(matrix_comp_reg_0_im); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1090 = comp_status == 4'h3 ? $signed(_GEN_578) : $signed(matrix_comp_reg_0_re); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1091 = comp_status == 4'h3 ? $signed(_GEN_611) : $signed(matrix_comp_reg_1_im); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1092 = comp_status == 4'h3 ? $signed(_GEN_612) : $signed(matrix_comp_reg_1_re); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1093 = comp_status == 4'h3 ? $signed(_GEN_645) : $signed(matrix_comp_reg_2_im); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1094 = comp_status == 4'h3 ? $signed(_GEN_646) : $signed(matrix_comp_reg_2_re); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1095 = comp_status == 4'h3 ? $signed(_GEN_679) : $signed(matrix_comp_reg_3_im); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1096 = comp_status == 4'h3 ? $signed(_GEN_680) : $signed(matrix_comp_reg_3_re); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1097 = comp_status == 4'h3 ? $signed(_GEN_713) : $signed(matrix_comp_reg_4_im); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1098 = comp_status == 4'h3 ? $signed(_GEN_714) : $signed(matrix_comp_reg_4_re); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1099 = comp_status == 4'h3 ? $signed(_GEN_747) : $signed(matrix_comp_reg_5_im); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1100 = comp_status == 4'h3 ? $signed(_GEN_748) : $signed(matrix_comp_reg_5_re); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1101 = comp_status == 4'h3 ? $signed(_GEN_781) : $signed(matrix_comp_reg_6_im); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1102 = comp_status == 4'h3 ? $signed(_GEN_782) : $signed(matrix_comp_reg_6_re); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1103 = comp_status == 4'h3 ? $signed(_GEN_815) : $signed(matrix_comp_reg_7_im); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1104 = comp_status == 4'h3 ? $signed(_GEN_816) : $signed(matrix_comp_reg_7_re); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1105 = comp_status == 4'h3 ? $signed(_GEN_849) : $signed(matrix_comp_reg_8_im); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1106 = comp_status == 4'h3 ? $signed(_GEN_850) : $signed(matrix_comp_reg_8_re); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1107 = comp_status == 4'h3 ? $signed(_GEN_883) : $signed(matrix_comp_reg_9_im); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1108 = comp_status == 4'h3 ? $signed(_GEN_884) : $signed(matrix_comp_reg_9_re); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1109 = comp_status == 4'h3 ? $signed(_GEN_917) : $signed(matrix_comp_reg_10_im); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1110 = comp_status == 4'h3 ? $signed(_GEN_918) : $signed(matrix_comp_reg_10_re); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1111 = comp_status == 4'h3 ? $signed(_GEN_951) : $signed(matrix_comp_reg_11_im); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1112 = comp_status == 4'h3 ? $signed(_GEN_952) : $signed(matrix_comp_reg_11_re); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1113 = comp_status == 4'h3 ? $signed(_GEN_985) : $signed(matrix_comp_reg_12_im); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1114 = comp_status == 4'h3 ? $signed(_GEN_986) : $signed(matrix_comp_reg_12_re); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1115 = comp_status == 4'h3 ? $signed(_GEN_1019) : $signed(matrix_comp_reg_13_im); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1116 = comp_status == 4'h3 ? $signed(_GEN_1020) : $signed(matrix_comp_reg_13_re); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1117 = comp_status == 4'h3 ? $signed(_GEN_1053) : $signed(matrix_comp_reg_14_im); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1118 = comp_status == 4'h3 ? $signed(_GEN_1054) : $signed(matrix_comp_reg_14_re); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1119 = comp_status == 4'h3 ? $signed(_GEN_1087) : $signed(matrix_comp_reg_15_im); // @[Cholesky_V1.scala 172:37 127:42]
  wire [63:0] _GEN_1120 = comp_status == 4'h3 ? $signed(_GEN_1088) : $signed(matrix_comp_reg_15_re); // @[Cholesky_V1.scala 172:37 127:42]
  wire [31:0] _GEN_1121 = comp_status == 4'h3 ? _point_index_T_1 : point_index; // @[Cholesky_V1.scala 172:37 181:19 128:34]
  wire [3:0] _GEN_1122 = comp_status == 4'h3 ? 4'h1 : comp_status; // @[Cholesky_V1.scala 172:37 182:19 129:34]
  wire [3:0] _GEN_1124 = comp_status == 4'h2 ? _GEN_544 : _GEN_1122; // @[Cholesky_V1.scala 166:37]
  wire [31:0] _GEN_1157 = comp_status == 4'h2 ? point_index : _GEN_1121; // @[Cholesky_V1.scala 128:34 166:37]
  cholesky_comp_unit cholesky_comp_unit ( // @[Cholesky_V1.scala 131:54]
    .clock(cholesky_comp_unit_clock),
    .reset(cholesky_comp_unit_reset),
    .io_reset(cholesky_comp_unit_io_reset),
    .io_ready(cholesky_comp_unit_io_ready),
    .io_matrixIn_0_re(cholesky_comp_unit_io_matrixIn_0_re),
    .io_matrixIn_0_im(cholesky_comp_unit_io_matrixIn_0_im),
    .io_matrixIn_1_re(cholesky_comp_unit_io_matrixIn_1_re),
    .io_matrixIn_1_im(cholesky_comp_unit_io_matrixIn_1_im),
    .io_matrixIn_2_re(cholesky_comp_unit_io_matrixIn_2_re),
    .io_matrixIn_2_im(cholesky_comp_unit_io_matrixIn_2_im),
    .io_matrixIn_3_re(cholesky_comp_unit_io_matrixIn_3_re),
    .io_matrixIn_3_im(cholesky_comp_unit_io_matrixIn_3_im),
    .io_matrixIn_4_re(cholesky_comp_unit_io_matrixIn_4_re),
    .io_matrixIn_4_im(cholesky_comp_unit_io_matrixIn_4_im),
    .io_matrixIn_5_re(cholesky_comp_unit_io_matrixIn_5_re),
    .io_matrixIn_5_im(cholesky_comp_unit_io_matrixIn_5_im),
    .io_matrixIn_6_re(cholesky_comp_unit_io_matrixIn_6_re),
    .io_matrixIn_6_im(cholesky_comp_unit_io_matrixIn_6_im),
    .io_matrixIn_7_re(cholesky_comp_unit_io_matrixIn_7_re),
    .io_matrixIn_7_im(cholesky_comp_unit_io_matrixIn_7_im),
    .io_matrixIn_8_re(cholesky_comp_unit_io_matrixIn_8_re),
    .io_matrixIn_8_im(cholesky_comp_unit_io_matrixIn_8_im),
    .io_matrixIn_9_re(cholesky_comp_unit_io_matrixIn_9_re),
    .io_matrixIn_9_im(cholesky_comp_unit_io_matrixIn_9_im),
    .io_matrixIn_10_re(cholesky_comp_unit_io_matrixIn_10_re),
    .io_matrixIn_10_im(cholesky_comp_unit_io_matrixIn_10_im),
    .io_matrixIn_11_re(cholesky_comp_unit_io_matrixIn_11_re),
    .io_matrixIn_11_im(cholesky_comp_unit_io_matrixIn_11_im),
    .io_matrixIn_12_re(cholesky_comp_unit_io_matrixIn_12_re),
    .io_matrixIn_12_im(cholesky_comp_unit_io_matrixIn_12_im),
    .io_matrixIn_13_re(cholesky_comp_unit_io_matrixIn_13_re),
    .io_matrixIn_13_im(cholesky_comp_unit_io_matrixIn_13_im),
    .io_matrixIn_14_re(cholesky_comp_unit_io_matrixIn_14_re),
    .io_matrixIn_14_im(cholesky_comp_unit_io_matrixIn_14_im),
    .io_matrixIn_15_re(cholesky_comp_unit_io_matrixIn_15_re),
    .io_matrixIn_15_im(cholesky_comp_unit_io_matrixIn_15_im),
    .io_matrixOut_0_re(cholesky_comp_unit_io_matrixOut_0_re),
    .io_matrixOut_0_im(cholesky_comp_unit_io_matrixOut_0_im),
    .io_matrixOut_1_re(cholesky_comp_unit_io_matrixOut_1_re),
    .io_matrixOut_1_im(cholesky_comp_unit_io_matrixOut_1_im),
    .io_matrixOut_2_re(cholesky_comp_unit_io_matrixOut_2_re),
    .io_matrixOut_2_im(cholesky_comp_unit_io_matrixOut_2_im),
    .io_matrixOut_3_re(cholesky_comp_unit_io_matrixOut_3_re),
    .io_matrixOut_3_im(cholesky_comp_unit_io_matrixOut_3_im),
    .io_matrixOut_4_re(cholesky_comp_unit_io_matrixOut_4_re),
    .io_matrixOut_4_im(cholesky_comp_unit_io_matrixOut_4_im),
    .io_matrixOut_5_re(cholesky_comp_unit_io_matrixOut_5_re),
    .io_matrixOut_5_im(cholesky_comp_unit_io_matrixOut_5_im),
    .io_matrixOut_6_re(cholesky_comp_unit_io_matrixOut_6_re),
    .io_matrixOut_6_im(cholesky_comp_unit_io_matrixOut_6_im),
    .io_matrixOut_7_re(cholesky_comp_unit_io_matrixOut_7_re),
    .io_matrixOut_7_im(cholesky_comp_unit_io_matrixOut_7_im),
    .io_matrixOut_8_re(cholesky_comp_unit_io_matrixOut_8_re),
    .io_matrixOut_8_im(cholesky_comp_unit_io_matrixOut_8_im),
    .io_matrixOut_9_re(cholesky_comp_unit_io_matrixOut_9_re),
    .io_matrixOut_9_im(cholesky_comp_unit_io_matrixOut_9_im),
    .io_matrixOut_10_re(cholesky_comp_unit_io_matrixOut_10_re),
    .io_matrixOut_10_im(cholesky_comp_unit_io_matrixOut_10_im),
    .io_matrixOut_11_re(cholesky_comp_unit_io_matrixOut_11_re),
    .io_matrixOut_11_im(cholesky_comp_unit_io_matrixOut_11_im),
    .io_matrixOut_12_re(cholesky_comp_unit_io_matrixOut_12_re),
    .io_matrixOut_12_im(cholesky_comp_unit_io_matrixOut_12_im),
    .io_matrixOut_13_re(cholesky_comp_unit_io_matrixOut_13_re),
    .io_matrixOut_13_im(cholesky_comp_unit_io_matrixOut_13_im),
    .io_matrixOut_14_re(cholesky_comp_unit_io_matrixOut_14_re),
    .io_matrixOut_14_im(cholesky_comp_unit_io_matrixOut_14_im),
    .io_matrixOut_15_re(cholesky_comp_unit_io_matrixOut_15_re),
    .io_matrixOut_15_im(cholesky_comp_unit_io_matrixOut_15_im),
    .io_valid(cholesky_comp_unit_io_valid)
  );
  assign io_matrixOut_0_re = matrix_comp_reg_0_re; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_0_im = matrix_comp_reg_0_im; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_1_re = matrix_comp_reg_4_re; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_1_im = matrix_comp_reg_4_im; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_2_re = matrix_comp_reg_5_re; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_2_im = matrix_comp_reg_5_im; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_3_re = matrix_comp_reg_8_re; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_3_im = matrix_comp_reg_8_im; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_4_re = matrix_comp_reg_9_re; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_4_im = matrix_comp_reg_9_im; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_5_re = matrix_comp_reg_10_re; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_5_im = matrix_comp_reg_10_im; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_6_re = matrix_comp_reg_12_re; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_6_im = matrix_comp_reg_12_im; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_7_re = matrix_comp_reg_13_re; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_7_im = matrix_comp_reg_13_im; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_8_re = matrix_comp_reg_14_re; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_8_im = matrix_comp_reg_14_im; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_9_re = matrix_comp_reg_15_re; // @[Cholesky_V1.scala 195:27]
  assign io_matrixOut_9_im = matrix_comp_reg_15_im; // @[Cholesky_V1.scala 195:27]
  assign io_valid = point_index >= 32'h4; // @[Cholesky_V1.scala 186:20]
  assign cholesky_comp_unit_clock = clock;
  assign cholesky_comp_unit_reset = reset;
  assign cholesky_comp_unit_io_reset = io_reset; // @[Cholesky_V1.scala 132:31]
  assign cholesky_comp_unit_io_ready = comp_status == 4'h1; // @[Cholesky_V1.scala 151:22]
  assign cholesky_comp_unit_io_matrixIn_0_re = 32'h0 < _T_2 & 32'h0 < _T_2 ? $signed(_GEN_31) : $signed(64'sh0); // @[Cholesky_V1.scala 157:76 158:55 161:58]
  assign cholesky_comp_unit_io_matrixIn_0_im = 4'hf == _cholesky_comp_unit_io_matrixIn_0_T_6[3:0] ? $signed(
    matrix_comp_reg_15_im) : $signed(_GEN_14); // @[Cholesky_V1.scala 158:{55,55}]
  assign cholesky_comp_unit_io_matrixIn_1_re = 32'h0 < _T_2 & 32'h1 < _T_2 ? $signed(_GEN_65) : $signed(64'sh0); // @[Cholesky_V1.scala 157:76 158:55 161:58]
  assign cholesky_comp_unit_io_matrixIn_1_im = 4'hf == _cholesky_comp_unit_io_matrixIn_1_T_6[3:0] ? $signed(
    matrix_comp_reg_15_im) : $signed(_GEN_48); // @[Cholesky_V1.scala 158:{55,55}]
  assign cholesky_comp_unit_io_matrixIn_2_re = 32'h0 < _T_2 & 32'h2 < _T_2 ? $signed(_GEN_99) : $signed(64'sh0); // @[Cholesky_V1.scala 157:76 158:55 161:58]
  assign cholesky_comp_unit_io_matrixIn_2_im = 4'hf == _cholesky_comp_unit_io_matrixIn_2_T_6[3:0] ? $signed(
    matrix_comp_reg_15_im) : $signed(_GEN_82); // @[Cholesky_V1.scala 158:{55,55}]
  assign cholesky_comp_unit_io_matrixIn_3_re = 32'h0 < _T_2 & 32'h3 < _T_2 ? $signed(_GEN_133) : $signed(64'sh0); // @[Cholesky_V1.scala 157:76 158:55 161:58]
  assign cholesky_comp_unit_io_matrixIn_3_im = 4'hf == _cholesky_comp_unit_io_matrixIn_3_T_6[3:0] ? $signed(
    matrix_comp_reg_15_im) : $signed(_GEN_116); // @[Cholesky_V1.scala 158:{55,55}]
  assign cholesky_comp_unit_io_matrixIn_4_re = 32'h1 < _T_2 & 32'h0 < _T_2 ? $signed(_GEN_167) : $signed(64'sh0); // @[Cholesky_V1.scala 157:76 158:55 161:58]
  assign cholesky_comp_unit_io_matrixIn_4_im = 4'hf == _cholesky_comp_unit_io_matrixIn_4_T_6[3:0] ? $signed(
    matrix_comp_reg_15_im) : $signed(_GEN_150); // @[Cholesky_V1.scala 158:{55,55}]
  assign cholesky_comp_unit_io_matrixIn_5_re = 32'h1 < _T_2 & 32'h1 < _T_2 ? $signed(_GEN_201) : $signed(64'sh0); // @[Cholesky_V1.scala 157:76 158:55 161:58]
  assign cholesky_comp_unit_io_matrixIn_5_im = 4'hf == _cholesky_comp_unit_io_matrixIn_5_T_6[3:0] ? $signed(
    matrix_comp_reg_15_im) : $signed(_GEN_184); // @[Cholesky_V1.scala 158:{55,55}]
  assign cholesky_comp_unit_io_matrixIn_6_re = 32'h1 < _T_2 & 32'h2 < _T_2 ? $signed(_GEN_235) : $signed(64'sh0); // @[Cholesky_V1.scala 157:76 158:55 161:58]
  assign cholesky_comp_unit_io_matrixIn_6_im = 4'hf == _cholesky_comp_unit_io_matrixIn_6_T_6[3:0] ? $signed(
    matrix_comp_reg_15_im) : $signed(_GEN_218); // @[Cholesky_V1.scala 158:{55,55}]
  assign cholesky_comp_unit_io_matrixIn_7_re = 32'h1 < _T_2 & 32'h3 < _T_2 ? $signed(_GEN_269) : $signed(64'sh0); // @[Cholesky_V1.scala 157:76 158:55 161:58]
  assign cholesky_comp_unit_io_matrixIn_7_im = 4'hf == _cholesky_comp_unit_io_matrixIn_7_T_6[3:0] ? $signed(
    matrix_comp_reg_15_im) : $signed(_GEN_252); // @[Cholesky_V1.scala 158:{55,55}]
  assign cholesky_comp_unit_io_matrixIn_8_re = 32'h2 < _T_2 & 32'h0 < _T_2 ? $signed(_GEN_303) : $signed(64'sh0); // @[Cholesky_V1.scala 157:76 158:55 161:58]
  assign cholesky_comp_unit_io_matrixIn_8_im = 4'hf == _cholesky_comp_unit_io_matrixIn_8_T_6[3:0] ? $signed(
    matrix_comp_reg_15_im) : $signed(_GEN_286); // @[Cholesky_V1.scala 158:{55,55}]
  assign cholesky_comp_unit_io_matrixIn_9_re = 32'h2 < _T_2 & 32'h1 < _T_2 ? $signed(_GEN_337) : $signed(64'sh0); // @[Cholesky_V1.scala 157:76 158:55 161:58]
  assign cholesky_comp_unit_io_matrixIn_9_im = 4'hf == _cholesky_comp_unit_io_matrixIn_9_T_6[3:0] ? $signed(
    matrix_comp_reg_15_im) : $signed(_GEN_320); // @[Cholesky_V1.scala 158:{55,55}]
  assign cholesky_comp_unit_io_matrixIn_10_re = 32'h2 < _T_2 & 32'h2 < _T_2 ? $signed(_GEN_371) : $signed(64'sh0); // @[Cholesky_V1.scala 157:76 158:55 161:58]
  assign cholesky_comp_unit_io_matrixIn_10_im = 4'hf == _cholesky_comp_unit_io_matrixIn_10_T_6[3:0] ? $signed(
    matrix_comp_reg_15_im) : $signed(_GEN_354); // @[Cholesky_V1.scala 158:{55,55}]
  assign cholesky_comp_unit_io_matrixIn_11_re = 32'h2 < _T_2 & 32'h3 < _T_2 ? $signed(_GEN_405) : $signed(64'sh0); // @[Cholesky_V1.scala 157:76 158:55 161:58]
  assign cholesky_comp_unit_io_matrixIn_11_im = 4'hf == _cholesky_comp_unit_io_matrixIn_11_T_6[3:0] ? $signed(
    matrix_comp_reg_15_im) : $signed(_GEN_388); // @[Cholesky_V1.scala 158:{55,55}]
  assign cholesky_comp_unit_io_matrixIn_12_re = 32'h3 < _T_2 & 32'h0 < _T_2 ? $signed(_GEN_439) : $signed(64'sh0); // @[Cholesky_V1.scala 157:76 158:55 161:58]
  assign cholesky_comp_unit_io_matrixIn_12_im = 4'hf == _cholesky_comp_unit_io_matrixIn_12_T_6[3:0] ? $signed(
    matrix_comp_reg_15_im) : $signed(_GEN_422); // @[Cholesky_V1.scala 158:{55,55}]
  assign cholesky_comp_unit_io_matrixIn_13_re = 32'h3 < _T_2 & 32'h1 < _T_2 ? $signed(_GEN_473) : $signed(64'sh0); // @[Cholesky_V1.scala 157:76 158:55 161:58]
  assign cholesky_comp_unit_io_matrixIn_13_im = 4'hf == _cholesky_comp_unit_io_matrixIn_13_T_6[3:0] ? $signed(
    matrix_comp_reg_15_im) : $signed(_GEN_456); // @[Cholesky_V1.scala 158:{55,55}]
  assign cholesky_comp_unit_io_matrixIn_14_re = 32'h3 < _T_2 & 32'h2 < _T_2 ? $signed(_GEN_507) : $signed(64'sh0); // @[Cholesky_V1.scala 157:76 158:55 161:58]
  assign cholesky_comp_unit_io_matrixIn_14_im = 4'hf == _cholesky_comp_unit_io_matrixIn_14_T_6[3:0] ? $signed(
    matrix_comp_reg_15_im) : $signed(_GEN_490); // @[Cholesky_V1.scala 158:{55,55}]
  assign cholesky_comp_unit_io_matrixIn_15_re = 32'h3 < _T_2 & 32'h3 < _T_2 ? $signed(_GEN_541) : $signed(64'sh0); // @[Cholesky_V1.scala 157:76 158:55 161:58]
  assign cholesky_comp_unit_io_matrixIn_15_im = 4'hf == _cholesky_comp_unit_io_matrixIn_15_T_6[3:0] ? $signed(
    matrix_comp_reg_15_im) : $signed(_GEN_524); // @[Cholesky_V1.scala 158:{55,55}]
  always @(posedge clock) begin
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_0_re <= 64'sh0; // @[Cholesky_V1.scala 139:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_0_re <= io_matrixIn_0_re; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_0_re <= _GEN_1090;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_0_im <= 64'sh0; // @[Cholesky_V1.scala 140:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_0_im <= io_matrixIn_0_im; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_0_im <= _GEN_1089;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_1_re <= 64'sh0; // @[Cholesky_V1.scala 139:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_1_re <= io_matrixIn_1_re; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_1_re <= _GEN_1092;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_1_im <= 64'sh0; // @[Cholesky_V1.scala 140:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_1_im <= io_matrixIn_1_im; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_1_im <= _GEN_1091;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_2_re <= 64'sh0; // @[Cholesky_V1.scala 139:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_2_re <= io_matrixIn_2_re; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_2_re <= _GEN_1094;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_2_im <= 64'sh0; // @[Cholesky_V1.scala 140:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_2_im <= io_matrixIn_2_im; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_2_im <= _GEN_1093;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_3_re <= 64'sh0; // @[Cholesky_V1.scala 139:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_3_re <= io_matrixIn_3_re; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_3_re <= _GEN_1096;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_3_im <= 64'sh0; // @[Cholesky_V1.scala 140:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_3_im <= io_matrixIn_3_im; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_3_im <= _GEN_1095;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_4_re <= 64'sh0; // @[Cholesky_V1.scala 139:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_4_re <= io_matrixIn_4_re; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_4_re <= _GEN_1098;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_4_im <= 64'sh0; // @[Cholesky_V1.scala 140:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_4_im <= io_matrixIn_4_im; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_4_im <= _GEN_1097;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_5_re <= 64'sh0; // @[Cholesky_V1.scala 139:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_5_re <= io_matrixIn_5_re; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_5_re <= _GEN_1100;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_5_im <= 64'sh0; // @[Cholesky_V1.scala 140:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_5_im <= io_matrixIn_5_im; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_5_im <= _GEN_1099;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_6_re <= 64'sh0; // @[Cholesky_V1.scala 139:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_6_re <= io_matrixIn_6_re; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_6_re <= _GEN_1102;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_6_im <= 64'sh0; // @[Cholesky_V1.scala 140:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_6_im <= io_matrixIn_6_im; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_6_im <= _GEN_1101;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_7_re <= 64'sh0; // @[Cholesky_V1.scala 139:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_7_re <= io_matrixIn_7_re; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_7_re <= _GEN_1104;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_7_im <= 64'sh0; // @[Cholesky_V1.scala 140:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_7_im <= io_matrixIn_7_im; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_7_im <= _GEN_1103;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_8_re <= 64'sh0; // @[Cholesky_V1.scala 139:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_8_re <= io_matrixIn_8_re; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_8_re <= _GEN_1106;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_8_im <= 64'sh0; // @[Cholesky_V1.scala 140:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_8_im <= io_matrixIn_8_im; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_8_im <= _GEN_1105;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_9_re <= 64'sh0; // @[Cholesky_V1.scala 139:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_9_re <= io_matrixIn_9_re; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_9_re <= _GEN_1108;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_9_im <= 64'sh0; // @[Cholesky_V1.scala 140:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_9_im <= io_matrixIn_9_im; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_9_im <= _GEN_1107;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_10_re <= 64'sh0; // @[Cholesky_V1.scala 139:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_10_re <= io_matrixIn_10_re; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_10_re <= _GEN_1110;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_10_im <= 64'sh0; // @[Cholesky_V1.scala 140:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_10_im <= io_matrixIn_10_im; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_10_im <= _GEN_1109;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_11_re <= 64'sh0; // @[Cholesky_V1.scala 139:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_11_re <= io_matrixIn_11_re; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_11_re <= _GEN_1112;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_11_im <= 64'sh0; // @[Cholesky_V1.scala 140:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_11_im <= io_matrixIn_11_im; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_11_im <= _GEN_1111;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_12_re <= 64'sh0; // @[Cholesky_V1.scala 139:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_12_re <= io_matrixIn_12_re; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_12_re <= _GEN_1114;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_12_im <= 64'sh0; // @[Cholesky_V1.scala 140:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_12_im <= io_matrixIn_12_im; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_12_im <= _GEN_1113;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_13_re <= 64'sh0; // @[Cholesky_V1.scala 139:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_13_re <= io_matrixIn_13_re; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_13_re <= _GEN_1116;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_13_im <= 64'sh0; // @[Cholesky_V1.scala 140:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_13_im <= io_matrixIn_13_im; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_13_im <= _GEN_1115;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_14_re <= 64'sh0; // @[Cholesky_V1.scala 139:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_14_re <= io_matrixIn_14_re; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_14_re <= _GEN_1118;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_14_im <= 64'sh0; // @[Cholesky_V1.scala 140:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_14_im <= io_matrixIn_14_im; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_14_im <= _GEN_1117;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_15_re <= 64'sh0; // @[Cholesky_V1.scala 139:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_15_re <= io_matrixIn_15_re; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_15_re <= _GEN_1120;
      end
    end
    if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      matrix_comp_reg_15_im <= 64'sh0; // @[Cholesky_V1.scala 140:29]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      matrix_comp_reg_15_im <= io_matrixIn_15_im; // @[Cholesky_V1.scala 146:21]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      if (!(comp_status == 4'h2)) begin // @[Cholesky_V1.scala 166:37]
        matrix_comp_reg_15_im <= _GEN_1119;
      end
    end
    if (reset) begin // @[Cholesky_V1.scala 128:34]
      point_index <= 32'h0; // @[Cholesky_V1.scala 128:34]
    end else if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      point_index <= 32'h0; // @[Cholesky_V1.scala 142:17]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      point_index <= 32'h0; // @[Cholesky_V1.scala 147:17]
    end else if (!(comp_status == 4'h1)) begin // @[Cholesky_V1.scala 151:31]
      point_index <= _GEN_1157;
    end
    if (reset) begin // @[Cholesky_V1.scala 129:34]
      comp_status <= 4'h0; // @[Cholesky_V1.scala 129:34]
    end else if (io_reset) begin // @[Cholesky_V1.scala 136:18]
      comp_status <= 4'h0; // @[Cholesky_V1.scala 143:17]
    end else if (io_ready) begin // @[Cholesky_V1.scala 144:24]
      comp_status <= 4'h1; // @[Cholesky_V1.scala 148:17]
    end else if (comp_status == 4'h1) begin // @[Cholesky_V1.scala 151:31]
      comp_status <= 4'h2; // @[Cholesky_V1.scala 165:19]
    end else begin
      comp_status <= _GEN_1124;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  matrix_comp_reg_0_re = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  matrix_comp_reg_0_im = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  matrix_comp_reg_1_re = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  matrix_comp_reg_1_im = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  matrix_comp_reg_2_re = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  matrix_comp_reg_2_im = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  matrix_comp_reg_3_re = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  matrix_comp_reg_3_im = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  matrix_comp_reg_4_re = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  matrix_comp_reg_4_im = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  matrix_comp_reg_5_re = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  matrix_comp_reg_5_im = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  matrix_comp_reg_6_re = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  matrix_comp_reg_6_im = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  matrix_comp_reg_7_re = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  matrix_comp_reg_7_im = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  matrix_comp_reg_8_re = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  matrix_comp_reg_8_im = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  matrix_comp_reg_9_re = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  matrix_comp_reg_9_im = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  matrix_comp_reg_10_re = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  matrix_comp_reg_10_im = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  matrix_comp_reg_11_re = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  matrix_comp_reg_11_im = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  matrix_comp_reg_12_re = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  matrix_comp_reg_12_im = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  matrix_comp_reg_13_re = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  matrix_comp_reg_13_im = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  matrix_comp_reg_14_re = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  matrix_comp_reg_14_im = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  matrix_comp_reg_15_re = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  matrix_comp_reg_15_im = _RAND_31[63:0];
  _RAND_32 = {1{`RANDOM}};
  point_index = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  comp_status = _RAND_33[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_FixedPoint(
  input         clock,
  input         io_reset,
  input  [63:0] io_in_x,
  input  [63:0] io_in_y,
  output [63:0] io_out_pe,
  output [63:0] io_out_x,
  output [63:0] io_out_y
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] pe_reg; // @[Matrix_FixedPoint_Mul.scala 29:31]
  reg [63:0] x_reg; // @[Matrix_FixedPoint_Mul.scala 30:30]
  reg [63:0] y_reg; // @[Matrix_FixedPoint_Mul.scala 31:30]
  wire [127:0] _pe_reg_T = $signed(io_in_x) * $signed(io_in_y); // @[Matrix_FixedPoint_Mul.scala 40:32]
  wire [95:0] _GEN_3 = {$signed(pe_reg), 32'h0}; // @[Matrix_FixedPoint_Mul.scala 40:22]
  wire [127:0] _GEN_4 = {{32{_GEN_3[95]}},_GEN_3}; // @[Matrix_FixedPoint_Mul.scala 40:22]
  wire [127:0] _pe_reg_T_3 = $signed(_GEN_4) + $signed(_pe_reg_T); // @[Matrix_FixedPoint_Mul.scala 40:22]
  wire [127:0] _GEN_0 = io_reset ? $signed(128'sh0) : $signed(_pe_reg_T_3); // @[Matrix_FixedPoint_Mul.scala 33:18 35:12 40:12]
  wire [95:0] _GEN_5 = _GEN_0[127:32];
  assign io_out_pe = pe_reg; // @[Matrix_FixedPoint_Mul.scala 47:13]
  assign io_out_x = x_reg; // @[Matrix_FixedPoint_Mul.scala 48:12]
  assign io_out_y = y_reg; // @[Matrix_FixedPoint_Mul.scala 49:12]
  always @(posedge clock) begin
    pe_reg <= _GEN_5[63:0];
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 33:18]
      x_reg <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 36:11]
    end else begin
      x_reg <= io_in_x; // @[Matrix_FixedPoint_Mul.scala 42:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 33:18]
      y_reg <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 37:11]
    end else begin
      y_reg <= io_in_y; // @[Matrix_FixedPoint_Mul.scala 43:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pe_reg = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  x_reg = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  y_reg = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module matrix_fixedPoint_mul(
  input         clock,
  input         io_reset,
  input         io_ready,
  input  [63:0] io_matrixA_0,
  input  [63:0] io_matrixA_4,
  input  [63:0] io_matrixA_5,
  input  [63:0] io_matrixA_8,
  input  [63:0] io_matrixA_9,
  input  [63:0] io_matrixA_10,
  input  [63:0] io_matrixA_12,
  input  [63:0] io_matrixA_13,
  input  [63:0] io_matrixA_14,
  input  [63:0] io_matrixA_15,
  input  [63:0] io_matrixB_0,
  input  [63:0] io_matrixB_4,
  input  [63:0] io_matrixB_5,
  input  [63:0] io_matrixB_8,
  input  [63:0] io_matrixB_9,
  input  [63:0] io_matrixB_10,
  input  [63:0] io_matrixB_12,
  input  [63:0] io_matrixB_13,
  input  [63:0] io_matrixB_14,
  input  [63:0] io_matrixB_15,
  output [63:0] io_matrixC_0,
  output [63:0] io_matrixC_4,
  output [63:0] io_matrixC_5,
  output [63:0] io_matrixC_8,
  output [63:0] io_matrixC_9,
  output [63:0] io_matrixC_10,
  output [63:0] io_matrixC_12,
  output [63:0] io_matrixC_13,
  output [63:0] io_matrixC_14,
  output [63:0] io_matrixC_15,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire  PE_FixedPoint_clock; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_io_reset; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_io_in_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_io_in_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_io_out_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_io_out_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_1_clock; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_1_io_reset; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_1_io_in_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_1_io_in_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_1_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_1_io_out_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_1_io_out_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_2_clock; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_2_io_reset; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_2_io_in_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_2_io_in_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_2_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_2_io_out_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_2_io_out_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_3_clock; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_3_io_reset; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_3_io_in_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_3_io_in_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_3_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_3_io_out_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_3_io_out_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_4_clock; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_4_io_reset; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_4_io_in_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_4_io_in_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_4_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_4_io_out_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_4_io_out_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_5_clock; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_5_io_reset; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_5_io_in_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_5_io_in_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_5_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_5_io_out_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_5_io_out_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_6_clock; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_6_io_reset; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_6_io_in_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_6_io_in_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_6_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_6_io_out_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_6_io_out_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_7_clock; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_7_io_reset; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_7_io_in_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_7_io_in_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_7_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_7_io_out_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_7_io_out_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_8_clock; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_8_io_reset; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_8_io_in_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_8_io_in_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_8_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_8_io_out_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_8_io_out_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_9_clock; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_9_io_reset; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_9_io_in_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_9_io_in_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_9_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_9_io_out_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_9_io_out_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_10_clock; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_10_io_reset; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_10_io_in_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_10_io_in_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_10_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_10_io_out_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_10_io_out_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_11_clock; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_11_io_reset; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_11_io_in_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_11_io_in_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_11_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_11_io_out_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_11_io_out_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_12_clock; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_12_io_reset; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_12_io_in_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_12_io_in_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_12_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_12_io_out_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_12_io_out_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_13_clock; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_13_io_reset; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_13_io_in_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_13_io_in_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_13_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_13_io_out_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_13_io_out_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_14_clock; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_14_io_reset; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_14_io_in_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_14_io_in_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_14_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_14_io_out_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_14_io_out_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_15_clock; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire  PE_FixedPoint_15_io_reset; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_15_io_in_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_15_io_in_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_15_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_15_io_out_x; // @[Matrix_FixedPoint_Mul.scala 83:35]
  wire [63:0] PE_FixedPoint_15_io_out_y; // @[Matrix_FixedPoint_Mul.scala 83:35]
  reg [63:0] regsA_0; // @[Matrix_FixedPoint_Mul.scala 79:35]
  reg [63:0] regsA_4; // @[Matrix_FixedPoint_Mul.scala 79:35]
  reg [63:0] regsA_5; // @[Matrix_FixedPoint_Mul.scala 79:35]
  reg [63:0] regsA_8; // @[Matrix_FixedPoint_Mul.scala 79:35]
  reg [63:0] regsA_9; // @[Matrix_FixedPoint_Mul.scala 79:35]
  reg [63:0] regsA_10; // @[Matrix_FixedPoint_Mul.scala 79:35]
  reg [63:0] regsA_12; // @[Matrix_FixedPoint_Mul.scala 79:35]
  reg [63:0] regsA_13; // @[Matrix_FixedPoint_Mul.scala 79:35]
  reg [63:0] regsA_14; // @[Matrix_FixedPoint_Mul.scala 79:35]
  reg [63:0] regsA_15; // @[Matrix_FixedPoint_Mul.scala 79:35]
  reg [63:0] regsB_0; // @[Matrix_FixedPoint_Mul.scala 80:35]
  reg [63:0] regsB_4; // @[Matrix_FixedPoint_Mul.scala 80:35]
  reg [63:0] regsB_5; // @[Matrix_FixedPoint_Mul.scala 80:35]
  reg [63:0] regsB_8; // @[Matrix_FixedPoint_Mul.scala 80:35]
  reg [63:0] regsB_9; // @[Matrix_FixedPoint_Mul.scala 80:35]
  reg [63:0] regsB_10; // @[Matrix_FixedPoint_Mul.scala 80:35]
  reg [63:0] regsB_12; // @[Matrix_FixedPoint_Mul.scala 80:35]
  reg [63:0] regsB_13; // @[Matrix_FixedPoint_Mul.scala 80:35]
  reg [63:0] regsB_14; // @[Matrix_FixedPoint_Mul.scala 80:35]
  reg [63:0] regsB_15; // @[Matrix_FixedPoint_Mul.scala 80:35]
  reg [4:0] input_point; // @[Matrix_FixedPoint_Mul.scala 81:30]
  wire [4:0] _input_point_T_1 = input_point + 5'h1; // @[Matrix_FixedPoint_Mul.scala 110:32]
  wire  _T = input_point < 5'h7; // @[Matrix_FixedPoint_Mul.scala 137:20]
  wire [3:0] _T_1 = 1'h0 * 3'h7; // @[Matrix_FixedPoint_Mul.scala 140:44]
  wire [4:0] _GEN_301 = {{1'd0}, _T_1}; // @[Matrix_FixedPoint_Mul.scala 140:60]
  wire [4:0] _T_3 = _GEN_301 + input_point; // @[Matrix_FixedPoint_Mul.scala 140:60]
  wire [63:0] _GEN_69 = 5'h1 == _T_3 ? $signed(64'sh0) : $signed(regsA_0); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_70 = 5'h2 == _T_3 ? $signed(64'sh0) : $signed(_GEN_69); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_71 = 5'h3 == _T_3 ? $signed(64'sh0) : $signed(_GEN_70); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_72 = 5'h4 == _T_3 ? $signed(64'sh0) : $signed(_GEN_71); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_73 = 5'h5 == _T_3 ? $signed(64'sh0) : $signed(_GEN_72); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_74 = 5'h6 == _T_3 ? $signed(64'sh0) : $signed(_GEN_73); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_75 = 5'h7 == _T_3 ? $signed(64'sh0) : $signed(_GEN_74); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_76 = 5'h8 == _T_3 ? $signed(regsA_4) : $signed(_GEN_75); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_77 = 5'h9 == _T_3 ? $signed(regsA_5) : $signed(_GEN_76); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_78 = 5'ha == _T_3 ? $signed(64'sh0) : $signed(_GEN_77); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_79 = 5'hb == _T_3 ? $signed(64'sh0) : $signed(_GEN_78); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_80 = 5'hc == _T_3 ? $signed(64'sh0) : $signed(_GEN_79); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_81 = 5'hd == _T_3 ? $signed(64'sh0) : $signed(_GEN_80); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_82 = 5'he == _T_3 ? $signed(64'sh0) : $signed(_GEN_81); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_83 = 5'hf == _T_3 ? $signed(64'sh0) : $signed(_GEN_82); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_84 = 5'h10 == _T_3 ? $signed(regsA_8) : $signed(_GEN_83); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_85 = 5'h11 == _T_3 ? $signed(regsA_9) : $signed(_GEN_84); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_86 = 5'h12 == _T_3 ? $signed(regsA_10) : $signed(_GEN_85); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_87 = 5'h13 == _T_3 ? $signed(64'sh0) : $signed(_GEN_86); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_88 = 5'h14 == _T_3 ? $signed(64'sh0) : $signed(_GEN_87); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_89 = 5'h15 == _T_3 ? $signed(64'sh0) : $signed(_GEN_88); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_90 = 5'h16 == _T_3 ? $signed(64'sh0) : $signed(_GEN_89); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_91 = 5'h17 == _T_3 ? $signed(64'sh0) : $signed(_GEN_90); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_92 = 5'h18 == _T_3 ? $signed(regsA_12) : $signed(_GEN_91); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_93 = 5'h19 == _T_3 ? $signed(regsA_13) : $signed(_GEN_92); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_94 = 5'h1a == _T_3 ? $signed(regsA_14) : $signed(_GEN_93); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_95 = 5'h1b == _T_3 ? $signed(regsA_15) : $signed(_GEN_94); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [3:0] _T_4 = 1'h1 * 3'h7; // @[Matrix_FixedPoint_Mul.scala 140:44]
  wire [4:0] _GEN_302 = {{1'd0}, _T_4}; // @[Matrix_FixedPoint_Mul.scala 140:60]
  wire [4:0] _T_6 = _GEN_302 + input_point; // @[Matrix_FixedPoint_Mul.scala 140:60]
  wire [63:0] _GEN_97 = 5'h1 == _T_6 ? $signed(64'sh0) : $signed(regsA_0); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_98 = 5'h2 == _T_6 ? $signed(64'sh0) : $signed(_GEN_97); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_99 = 5'h3 == _T_6 ? $signed(64'sh0) : $signed(_GEN_98); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_100 = 5'h4 == _T_6 ? $signed(64'sh0) : $signed(_GEN_99); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_101 = 5'h5 == _T_6 ? $signed(64'sh0) : $signed(_GEN_100); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_102 = 5'h6 == _T_6 ? $signed(64'sh0) : $signed(_GEN_101); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_103 = 5'h7 == _T_6 ? $signed(64'sh0) : $signed(_GEN_102); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_104 = 5'h8 == _T_6 ? $signed(regsA_4) : $signed(_GEN_103); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_105 = 5'h9 == _T_6 ? $signed(regsA_5) : $signed(_GEN_104); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_106 = 5'ha == _T_6 ? $signed(64'sh0) : $signed(_GEN_105); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_107 = 5'hb == _T_6 ? $signed(64'sh0) : $signed(_GEN_106); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_108 = 5'hc == _T_6 ? $signed(64'sh0) : $signed(_GEN_107); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_109 = 5'hd == _T_6 ? $signed(64'sh0) : $signed(_GEN_108); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_110 = 5'he == _T_6 ? $signed(64'sh0) : $signed(_GEN_109); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_111 = 5'hf == _T_6 ? $signed(64'sh0) : $signed(_GEN_110); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_112 = 5'h10 == _T_6 ? $signed(regsA_8) : $signed(_GEN_111); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_113 = 5'h11 == _T_6 ? $signed(regsA_9) : $signed(_GEN_112); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_114 = 5'h12 == _T_6 ? $signed(regsA_10) : $signed(_GEN_113); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_115 = 5'h13 == _T_6 ? $signed(64'sh0) : $signed(_GEN_114); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_116 = 5'h14 == _T_6 ? $signed(64'sh0) : $signed(_GEN_115); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_117 = 5'h15 == _T_6 ? $signed(64'sh0) : $signed(_GEN_116); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_118 = 5'h16 == _T_6 ? $signed(64'sh0) : $signed(_GEN_117); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_119 = 5'h17 == _T_6 ? $signed(64'sh0) : $signed(_GEN_118); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_120 = 5'h18 == _T_6 ? $signed(regsA_12) : $signed(_GEN_119); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_121 = 5'h19 == _T_6 ? $signed(regsA_13) : $signed(_GEN_120); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_122 = 5'h1a == _T_6 ? $signed(regsA_14) : $signed(_GEN_121); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_123 = 5'h1b == _T_6 ? $signed(regsA_15) : $signed(_GEN_122); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [4:0] _T_7 = 2'h2 * 3'h7; // @[Matrix_FixedPoint_Mul.scala 140:44]
  wire [4:0] _T_9 = _T_7 + input_point; // @[Matrix_FixedPoint_Mul.scala 140:60]
  wire [63:0] _GEN_125 = 5'h1 == _T_9 ? $signed(64'sh0) : $signed(regsA_0); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_126 = 5'h2 == _T_9 ? $signed(64'sh0) : $signed(_GEN_125); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_127 = 5'h3 == _T_9 ? $signed(64'sh0) : $signed(_GEN_126); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_128 = 5'h4 == _T_9 ? $signed(64'sh0) : $signed(_GEN_127); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_129 = 5'h5 == _T_9 ? $signed(64'sh0) : $signed(_GEN_128); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_130 = 5'h6 == _T_9 ? $signed(64'sh0) : $signed(_GEN_129); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_131 = 5'h7 == _T_9 ? $signed(64'sh0) : $signed(_GEN_130); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_132 = 5'h8 == _T_9 ? $signed(regsA_4) : $signed(_GEN_131); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_133 = 5'h9 == _T_9 ? $signed(regsA_5) : $signed(_GEN_132); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_134 = 5'ha == _T_9 ? $signed(64'sh0) : $signed(_GEN_133); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_135 = 5'hb == _T_9 ? $signed(64'sh0) : $signed(_GEN_134); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_136 = 5'hc == _T_9 ? $signed(64'sh0) : $signed(_GEN_135); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_137 = 5'hd == _T_9 ? $signed(64'sh0) : $signed(_GEN_136); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_138 = 5'he == _T_9 ? $signed(64'sh0) : $signed(_GEN_137); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_139 = 5'hf == _T_9 ? $signed(64'sh0) : $signed(_GEN_138); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_140 = 5'h10 == _T_9 ? $signed(regsA_8) : $signed(_GEN_139); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_141 = 5'h11 == _T_9 ? $signed(regsA_9) : $signed(_GEN_140); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_142 = 5'h12 == _T_9 ? $signed(regsA_10) : $signed(_GEN_141); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_143 = 5'h13 == _T_9 ? $signed(64'sh0) : $signed(_GEN_142); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_144 = 5'h14 == _T_9 ? $signed(64'sh0) : $signed(_GEN_143); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_145 = 5'h15 == _T_9 ? $signed(64'sh0) : $signed(_GEN_144); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_146 = 5'h16 == _T_9 ? $signed(64'sh0) : $signed(_GEN_145); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_147 = 5'h17 == _T_9 ? $signed(64'sh0) : $signed(_GEN_146); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_148 = 5'h18 == _T_9 ? $signed(regsA_12) : $signed(_GEN_147); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_149 = 5'h19 == _T_9 ? $signed(regsA_13) : $signed(_GEN_148); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_150 = 5'h1a == _T_9 ? $signed(regsA_14) : $signed(_GEN_149); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_151 = 5'h1b == _T_9 ? $signed(regsA_15) : $signed(_GEN_150); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [4:0] _T_10 = 2'h3 * 3'h7; // @[Matrix_FixedPoint_Mul.scala 140:44]
  wire [4:0] _T_12 = _T_10 + input_point; // @[Matrix_FixedPoint_Mul.scala 140:60]
  wire [63:0] _GEN_153 = 5'h1 == _T_12 ? $signed(64'sh0) : $signed(regsA_0); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_154 = 5'h2 == _T_12 ? $signed(64'sh0) : $signed(_GEN_153); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_155 = 5'h3 == _T_12 ? $signed(64'sh0) : $signed(_GEN_154); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_156 = 5'h4 == _T_12 ? $signed(64'sh0) : $signed(_GEN_155); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_157 = 5'h5 == _T_12 ? $signed(64'sh0) : $signed(_GEN_156); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_158 = 5'h6 == _T_12 ? $signed(64'sh0) : $signed(_GEN_157); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_159 = 5'h7 == _T_12 ? $signed(64'sh0) : $signed(_GEN_158); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_160 = 5'h8 == _T_12 ? $signed(regsA_4) : $signed(_GEN_159); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_161 = 5'h9 == _T_12 ? $signed(regsA_5) : $signed(_GEN_160); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_162 = 5'ha == _T_12 ? $signed(64'sh0) : $signed(_GEN_161); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_163 = 5'hb == _T_12 ? $signed(64'sh0) : $signed(_GEN_162); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_164 = 5'hc == _T_12 ? $signed(64'sh0) : $signed(_GEN_163); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_165 = 5'hd == _T_12 ? $signed(64'sh0) : $signed(_GEN_164); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_166 = 5'he == _T_12 ? $signed(64'sh0) : $signed(_GEN_165); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_167 = 5'hf == _T_12 ? $signed(64'sh0) : $signed(_GEN_166); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_168 = 5'h10 == _T_12 ? $signed(regsA_8) : $signed(_GEN_167); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_169 = 5'h11 == _T_12 ? $signed(regsA_9) : $signed(_GEN_168); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_170 = 5'h12 == _T_12 ? $signed(regsA_10) : $signed(_GEN_169); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_171 = 5'h13 == _T_12 ? $signed(64'sh0) : $signed(_GEN_170); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_172 = 5'h14 == _T_12 ? $signed(64'sh0) : $signed(_GEN_171); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_173 = 5'h15 == _T_12 ? $signed(64'sh0) : $signed(_GEN_172); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_174 = 5'h16 == _T_12 ? $signed(64'sh0) : $signed(_GEN_173); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_175 = 5'h17 == _T_12 ? $signed(64'sh0) : $signed(_GEN_174); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_176 = 5'h18 == _T_12 ? $signed(regsA_12) : $signed(_GEN_175); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_177 = 5'h19 == _T_12 ? $signed(regsA_13) : $signed(_GEN_176); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_178 = 5'h1a == _T_12 ? $signed(regsA_14) : $signed(_GEN_177); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_179 = 5'h1b == _T_12 ? $signed(regsA_15) : $signed(_GEN_178); // @[Matrix_FixedPoint_Mul.scala 140:{27,27}]
  wire [63:0] _GEN_185 = 5'h1 == _T_3 ? $signed(regsB_4) : $signed(regsB_0); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_186 = 5'h2 == _T_3 ? $signed(regsB_8) : $signed(_GEN_185); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_187 = 5'h3 == _T_3 ? $signed(regsB_12) : $signed(_GEN_186); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_188 = 5'h4 == _T_3 ? $signed(64'sh0) : $signed(_GEN_187); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_189 = 5'h5 == _T_3 ? $signed(64'sh0) : $signed(_GEN_188); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_190 = 5'h6 == _T_3 ? $signed(64'sh0) : $signed(_GEN_189); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_191 = 5'h7 == _T_3 ? $signed(64'sh0) : $signed(_GEN_190); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_192 = 5'h8 == _T_3 ? $signed(64'sh0) : $signed(_GEN_191); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_193 = 5'h9 == _T_3 ? $signed(regsB_5) : $signed(_GEN_192); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_194 = 5'ha == _T_3 ? $signed(regsB_9) : $signed(_GEN_193); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_195 = 5'hb == _T_3 ? $signed(regsB_13) : $signed(_GEN_194); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_196 = 5'hc == _T_3 ? $signed(64'sh0) : $signed(_GEN_195); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_197 = 5'hd == _T_3 ? $signed(64'sh0) : $signed(_GEN_196); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_198 = 5'he == _T_3 ? $signed(64'sh0) : $signed(_GEN_197); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_199 = 5'hf == _T_3 ? $signed(64'sh0) : $signed(_GEN_198); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_200 = 5'h10 == _T_3 ? $signed(64'sh0) : $signed(_GEN_199); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_201 = 5'h11 == _T_3 ? $signed(64'sh0) : $signed(_GEN_200); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_202 = 5'h12 == _T_3 ? $signed(regsB_10) : $signed(_GEN_201); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_203 = 5'h13 == _T_3 ? $signed(regsB_14) : $signed(_GEN_202); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_204 = 5'h14 == _T_3 ? $signed(64'sh0) : $signed(_GEN_203); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_205 = 5'h15 == _T_3 ? $signed(64'sh0) : $signed(_GEN_204); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_206 = 5'h16 == _T_3 ? $signed(64'sh0) : $signed(_GEN_205); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_207 = 5'h17 == _T_3 ? $signed(64'sh0) : $signed(_GEN_206); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_208 = 5'h18 == _T_3 ? $signed(64'sh0) : $signed(_GEN_207); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_209 = 5'h19 == _T_3 ? $signed(64'sh0) : $signed(_GEN_208); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_210 = 5'h1a == _T_3 ? $signed(64'sh0) : $signed(_GEN_209); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_211 = 5'h1b == _T_3 ? $signed(regsB_15) : $signed(_GEN_210); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_213 = 5'h1 == _T_6 ? $signed(regsB_4) : $signed(regsB_0); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_214 = 5'h2 == _T_6 ? $signed(regsB_8) : $signed(_GEN_213); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_215 = 5'h3 == _T_6 ? $signed(regsB_12) : $signed(_GEN_214); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_216 = 5'h4 == _T_6 ? $signed(64'sh0) : $signed(_GEN_215); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_217 = 5'h5 == _T_6 ? $signed(64'sh0) : $signed(_GEN_216); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_218 = 5'h6 == _T_6 ? $signed(64'sh0) : $signed(_GEN_217); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_219 = 5'h7 == _T_6 ? $signed(64'sh0) : $signed(_GEN_218); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_220 = 5'h8 == _T_6 ? $signed(64'sh0) : $signed(_GEN_219); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_221 = 5'h9 == _T_6 ? $signed(regsB_5) : $signed(_GEN_220); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_222 = 5'ha == _T_6 ? $signed(regsB_9) : $signed(_GEN_221); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_223 = 5'hb == _T_6 ? $signed(regsB_13) : $signed(_GEN_222); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_224 = 5'hc == _T_6 ? $signed(64'sh0) : $signed(_GEN_223); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_225 = 5'hd == _T_6 ? $signed(64'sh0) : $signed(_GEN_224); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_226 = 5'he == _T_6 ? $signed(64'sh0) : $signed(_GEN_225); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_227 = 5'hf == _T_6 ? $signed(64'sh0) : $signed(_GEN_226); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_228 = 5'h10 == _T_6 ? $signed(64'sh0) : $signed(_GEN_227); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_229 = 5'h11 == _T_6 ? $signed(64'sh0) : $signed(_GEN_228); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_230 = 5'h12 == _T_6 ? $signed(regsB_10) : $signed(_GEN_229); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_231 = 5'h13 == _T_6 ? $signed(regsB_14) : $signed(_GEN_230); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_232 = 5'h14 == _T_6 ? $signed(64'sh0) : $signed(_GEN_231); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_233 = 5'h15 == _T_6 ? $signed(64'sh0) : $signed(_GEN_232); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_234 = 5'h16 == _T_6 ? $signed(64'sh0) : $signed(_GEN_233); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_235 = 5'h17 == _T_6 ? $signed(64'sh0) : $signed(_GEN_234); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_236 = 5'h18 == _T_6 ? $signed(64'sh0) : $signed(_GEN_235); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_237 = 5'h19 == _T_6 ? $signed(64'sh0) : $signed(_GEN_236); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_238 = 5'h1a == _T_6 ? $signed(64'sh0) : $signed(_GEN_237); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_239 = 5'h1b == _T_6 ? $signed(regsB_15) : $signed(_GEN_238); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_241 = 5'h1 == _T_9 ? $signed(regsB_4) : $signed(regsB_0); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_242 = 5'h2 == _T_9 ? $signed(regsB_8) : $signed(_GEN_241); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_243 = 5'h3 == _T_9 ? $signed(regsB_12) : $signed(_GEN_242); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_244 = 5'h4 == _T_9 ? $signed(64'sh0) : $signed(_GEN_243); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_245 = 5'h5 == _T_9 ? $signed(64'sh0) : $signed(_GEN_244); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_246 = 5'h6 == _T_9 ? $signed(64'sh0) : $signed(_GEN_245); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_247 = 5'h7 == _T_9 ? $signed(64'sh0) : $signed(_GEN_246); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_248 = 5'h8 == _T_9 ? $signed(64'sh0) : $signed(_GEN_247); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_249 = 5'h9 == _T_9 ? $signed(regsB_5) : $signed(_GEN_248); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_250 = 5'ha == _T_9 ? $signed(regsB_9) : $signed(_GEN_249); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_251 = 5'hb == _T_9 ? $signed(regsB_13) : $signed(_GEN_250); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_252 = 5'hc == _T_9 ? $signed(64'sh0) : $signed(_GEN_251); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_253 = 5'hd == _T_9 ? $signed(64'sh0) : $signed(_GEN_252); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_254 = 5'he == _T_9 ? $signed(64'sh0) : $signed(_GEN_253); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_255 = 5'hf == _T_9 ? $signed(64'sh0) : $signed(_GEN_254); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_256 = 5'h10 == _T_9 ? $signed(64'sh0) : $signed(_GEN_255); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_257 = 5'h11 == _T_9 ? $signed(64'sh0) : $signed(_GEN_256); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_258 = 5'h12 == _T_9 ? $signed(regsB_10) : $signed(_GEN_257); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_259 = 5'h13 == _T_9 ? $signed(regsB_14) : $signed(_GEN_258); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_260 = 5'h14 == _T_9 ? $signed(64'sh0) : $signed(_GEN_259); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_261 = 5'h15 == _T_9 ? $signed(64'sh0) : $signed(_GEN_260); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_262 = 5'h16 == _T_9 ? $signed(64'sh0) : $signed(_GEN_261); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_263 = 5'h17 == _T_9 ? $signed(64'sh0) : $signed(_GEN_262); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_264 = 5'h18 == _T_9 ? $signed(64'sh0) : $signed(_GEN_263); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_265 = 5'h19 == _T_9 ? $signed(64'sh0) : $signed(_GEN_264); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_266 = 5'h1a == _T_9 ? $signed(64'sh0) : $signed(_GEN_265); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_267 = 5'h1b == _T_9 ? $signed(regsB_15) : $signed(_GEN_266); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_269 = 5'h1 == _T_12 ? $signed(regsB_4) : $signed(regsB_0); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_270 = 5'h2 == _T_12 ? $signed(regsB_8) : $signed(_GEN_269); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_271 = 5'h3 == _T_12 ? $signed(regsB_12) : $signed(_GEN_270); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_272 = 5'h4 == _T_12 ? $signed(64'sh0) : $signed(_GEN_271); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_273 = 5'h5 == _T_12 ? $signed(64'sh0) : $signed(_GEN_272); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_274 = 5'h6 == _T_12 ? $signed(64'sh0) : $signed(_GEN_273); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_275 = 5'h7 == _T_12 ? $signed(64'sh0) : $signed(_GEN_274); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_276 = 5'h8 == _T_12 ? $signed(64'sh0) : $signed(_GEN_275); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_277 = 5'h9 == _T_12 ? $signed(regsB_5) : $signed(_GEN_276); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_278 = 5'ha == _T_12 ? $signed(regsB_9) : $signed(_GEN_277); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_279 = 5'hb == _T_12 ? $signed(regsB_13) : $signed(_GEN_278); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_280 = 5'hc == _T_12 ? $signed(64'sh0) : $signed(_GEN_279); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_281 = 5'hd == _T_12 ? $signed(64'sh0) : $signed(_GEN_280); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_282 = 5'he == _T_12 ? $signed(64'sh0) : $signed(_GEN_281); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_283 = 5'hf == _T_12 ? $signed(64'sh0) : $signed(_GEN_282); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_284 = 5'h10 == _T_12 ? $signed(64'sh0) : $signed(_GEN_283); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_285 = 5'h11 == _T_12 ? $signed(64'sh0) : $signed(_GEN_284); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_286 = 5'h12 == _T_12 ? $signed(regsB_10) : $signed(_GEN_285); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_287 = 5'h13 == _T_12 ? $signed(regsB_14) : $signed(_GEN_286); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_288 = 5'h14 == _T_12 ? $signed(64'sh0) : $signed(_GEN_287); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_289 = 5'h15 == _T_12 ? $signed(64'sh0) : $signed(_GEN_288); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_290 = 5'h16 == _T_12 ? $signed(64'sh0) : $signed(_GEN_289); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_291 = 5'h17 == _T_12 ? $signed(64'sh0) : $signed(_GEN_290); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_292 = 5'h18 == _T_12 ? $signed(64'sh0) : $signed(_GEN_291); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_293 = 5'h19 == _T_12 ? $signed(64'sh0) : $signed(_GEN_292); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_294 = 5'h1a == _T_12 ? $signed(64'sh0) : $signed(_GEN_293); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  wire [63:0] _GEN_295 = 5'h1b == _T_12 ? $signed(regsB_15) : $signed(_GEN_294); // @[Matrix_FixedPoint_Mul.scala 152:{19,19}]
  PE_FixedPoint PE_FixedPoint ( // @[Matrix_FixedPoint_Mul.scala 83:35]
    .clock(PE_FixedPoint_clock),
    .io_reset(PE_FixedPoint_io_reset),
    .io_in_x(PE_FixedPoint_io_in_x),
    .io_in_y(PE_FixedPoint_io_in_y),
    .io_out_pe(PE_FixedPoint_io_out_pe),
    .io_out_x(PE_FixedPoint_io_out_x),
    .io_out_y(PE_FixedPoint_io_out_y)
  );
  PE_FixedPoint PE_FixedPoint_1 ( // @[Matrix_FixedPoint_Mul.scala 83:35]
    .clock(PE_FixedPoint_1_clock),
    .io_reset(PE_FixedPoint_1_io_reset),
    .io_in_x(PE_FixedPoint_1_io_in_x),
    .io_in_y(PE_FixedPoint_1_io_in_y),
    .io_out_pe(PE_FixedPoint_1_io_out_pe),
    .io_out_x(PE_FixedPoint_1_io_out_x),
    .io_out_y(PE_FixedPoint_1_io_out_y)
  );
  PE_FixedPoint PE_FixedPoint_2 ( // @[Matrix_FixedPoint_Mul.scala 83:35]
    .clock(PE_FixedPoint_2_clock),
    .io_reset(PE_FixedPoint_2_io_reset),
    .io_in_x(PE_FixedPoint_2_io_in_x),
    .io_in_y(PE_FixedPoint_2_io_in_y),
    .io_out_pe(PE_FixedPoint_2_io_out_pe),
    .io_out_x(PE_FixedPoint_2_io_out_x),
    .io_out_y(PE_FixedPoint_2_io_out_y)
  );
  PE_FixedPoint PE_FixedPoint_3 ( // @[Matrix_FixedPoint_Mul.scala 83:35]
    .clock(PE_FixedPoint_3_clock),
    .io_reset(PE_FixedPoint_3_io_reset),
    .io_in_x(PE_FixedPoint_3_io_in_x),
    .io_in_y(PE_FixedPoint_3_io_in_y),
    .io_out_pe(PE_FixedPoint_3_io_out_pe),
    .io_out_x(PE_FixedPoint_3_io_out_x),
    .io_out_y(PE_FixedPoint_3_io_out_y)
  );
  PE_FixedPoint PE_FixedPoint_4 ( // @[Matrix_FixedPoint_Mul.scala 83:35]
    .clock(PE_FixedPoint_4_clock),
    .io_reset(PE_FixedPoint_4_io_reset),
    .io_in_x(PE_FixedPoint_4_io_in_x),
    .io_in_y(PE_FixedPoint_4_io_in_y),
    .io_out_pe(PE_FixedPoint_4_io_out_pe),
    .io_out_x(PE_FixedPoint_4_io_out_x),
    .io_out_y(PE_FixedPoint_4_io_out_y)
  );
  PE_FixedPoint PE_FixedPoint_5 ( // @[Matrix_FixedPoint_Mul.scala 83:35]
    .clock(PE_FixedPoint_5_clock),
    .io_reset(PE_FixedPoint_5_io_reset),
    .io_in_x(PE_FixedPoint_5_io_in_x),
    .io_in_y(PE_FixedPoint_5_io_in_y),
    .io_out_pe(PE_FixedPoint_5_io_out_pe),
    .io_out_x(PE_FixedPoint_5_io_out_x),
    .io_out_y(PE_FixedPoint_5_io_out_y)
  );
  PE_FixedPoint PE_FixedPoint_6 ( // @[Matrix_FixedPoint_Mul.scala 83:35]
    .clock(PE_FixedPoint_6_clock),
    .io_reset(PE_FixedPoint_6_io_reset),
    .io_in_x(PE_FixedPoint_6_io_in_x),
    .io_in_y(PE_FixedPoint_6_io_in_y),
    .io_out_pe(PE_FixedPoint_6_io_out_pe),
    .io_out_x(PE_FixedPoint_6_io_out_x),
    .io_out_y(PE_FixedPoint_6_io_out_y)
  );
  PE_FixedPoint PE_FixedPoint_7 ( // @[Matrix_FixedPoint_Mul.scala 83:35]
    .clock(PE_FixedPoint_7_clock),
    .io_reset(PE_FixedPoint_7_io_reset),
    .io_in_x(PE_FixedPoint_7_io_in_x),
    .io_in_y(PE_FixedPoint_7_io_in_y),
    .io_out_pe(PE_FixedPoint_7_io_out_pe),
    .io_out_x(PE_FixedPoint_7_io_out_x),
    .io_out_y(PE_FixedPoint_7_io_out_y)
  );
  PE_FixedPoint PE_FixedPoint_8 ( // @[Matrix_FixedPoint_Mul.scala 83:35]
    .clock(PE_FixedPoint_8_clock),
    .io_reset(PE_FixedPoint_8_io_reset),
    .io_in_x(PE_FixedPoint_8_io_in_x),
    .io_in_y(PE_FixedPoint_8_io_in_y),
    .io_out_pe(PE_FixedPoint_8_io_out_pe),
    .io_out_x(PE_FixedPoint_8_io_out_x),
    .io_out_y(PE_FixedPoint_8_io_out_y)
  );
  PE_FixedPoint PE_FixedPoint_9 ( // @[Matrix_FixedPoint_Mul.scala 83:35]
    .clock(PE_FixedPoint_9_clock),
    .io_reset(PE_FixedPoint_9_io_reset),
    .io_in_x(PE_FixedPoint_9_io_in_x),
    .io_in_y(PE_FixedPoint_9_io_in_y),
    .io_out_pe(PE_FixedPoint_9_io_out_pe),
    .io_out_x(PE_FixedPoint_9_io_out_x),
    .io_out_y(PE_FixedPoint_9_io_out_y)
  );
  PE_FixedPoint PE_FixedPoint_10 ( // @[Matrix_FixedPoint_Mul.scala 83:35]
    .clock(PE_FixedPoint_10_clock),
    .io_reset(PE_FixedPoint_10_io_reset),
    .io_in_x(PE_FixedPoint_10_io_in_x),
    .io_in_y(PE_FixedPoint_10_io_in_y),
    .io_out_pe(PE_FixedPoint_10_io_out_pe),
    .io_out_x(PE_FixedPoint_10_io_out_x),
    .io_out_y(PE_FixedPoint_10_io_out_y)
  );
  PE_FixedPoint PE_FixedPoint_11 ( // @[Matrix_FixedPoint_Mul.scala 83:35]
    .clock(PE_FixedPoint_11_clock),
    .io_reset(PE_FixedPoint_11_io_reset),
    .io_in_x(PE_FixedPoint_11_io_in_x),
    .io_in_y(PE_FixedPoint_11_io_in_y),
    .io_out_pe(PE_FixedPoint_11_io_out_pe),
    .io_out_x(PE_FixedPoint_11_io_out_x),
    .io_out_y(PE_FixedPoint_11_io_out_y)
  );
  PE_FixedPoint PE_FixedPoint_12 ( // @[Matrix_FixedPoint_Mul.scala 83:35]
    .clock(PE_FixedPoint_12_clock),
    .io_reset(PE_FixedPoint_12_io_reset),
    .io_in_x(PE_FixedPoint_12_io_in_x),
    .io_in_y(PE_FixedPoint_12_io_in_y),
    .io_out_pe(PE_FixedPoint_12_io_out_pe),
    .io_out_x(PE_FixedPoint_12_io_out_x),
    .io_out_y(PE_FixedPoint_12_io_out_y)
  );
  PE_FixedPoint PE_FixedPoint_13 ( // @[Matrix_FixedPoint_Mul.scala 83:35]
    .clock(PE_FixedPoint_13_clock),
    .io_reset(PE_FixedPoint_13_io_reset),
    .io_in_x(PE_FixedPoint_13_io_in_x),
    .io_in_y(PE_FixedPoint_13_io_in_y),
    .io_out_pe(PE_FixedPoint_13_io_out_pe),
    .io_out_x(PE_FixedPoint_13_io_out_x),
    .io_out_y(PE_FixedPoint_13_io_out_y)
  );
  PE_FixedPoint PE_FixedPoint_14 ( // @[Matrix_FixedPoint_Mul.scala 83:35]
    .clock(PE_FixedPoint_14_clock),
    .io_reset(PE_FixedPoint_14_io_reset),
    .io_in_x(PE_FixedPoint_14_io_in_x),
    .io_in_y(PE_FixedPoint_14_io_in_y),
    .io_out_pe(PE_FixedPoint_14_io_out_pe),
    .io_out_x(PE_FixedPoint_14_io_out_x),
    .io_out_y(PE_FixedPoint_14_io_out_y)
  );
  PE_FixedPoint PE_FixedPoint_15 ( // @[Matrix_FixedPoint_Mul.scala 83:35]
    .clock(PE_FixedPoint_15_clock),
    .io_reset(PE_FixedPoint_15_io_reset),
    .io_in_x(PE_FixedPoint_15_io_in_x),
    .io_in_y(PE_FixedPoint_15_io_in_y),
    .io_out_pe(PE_FixedPoint_15_io_out_pe),
    .io_out_x(PE_FixedPoint_15_io_out_x),
    .io_out_y(PE_FixedPoint_15_io_out_y)
  );
  assign io_matrixC_0 = PE_FixedPoint_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 184:19]
  assign io_matrixC_4 = PE_FixedPoint_4_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 184:19]
  assign io_matrixC_5 = PE_FixedPoint_5_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 184:19]
  assign io_matrixC_8 = PE_FixedPoint_8_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 184:19]
  assign io_matrixC_9 = PE_FixedPoint_9_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 184:19]
  assign io_matrixC_10 = PE_FixedPoint_10_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 184:19]
  assign io_matrixC_12 = PE_FixedPoint_12_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 184:19]
  assign io_matrixC_13 = PE_FixedPoint_13_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 184:19]
  assign io_matrixC_14 = PE_FixedPoint_14_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 184:19]
  assign io_matrixC_15 = PE_FixedPoint_15_io_out_pe; // @[Matrix_FixedPoint_Mul.scala 184:19]
  assign io_valid = input_point >= 5'ha; // @[Matrix_FixedPoint_Mul.scala 177:20]
  assign PE_FixedPoint_clock = clock;
  assign PE_FixedPoint_io_reset = io_reset | io_ready; // @[Matrix_FixedPoint_Mul.scala 85:18 95:20]
  assign PE_FixedPoint_io_in_x = input_point < 5'h7 ? $signed(_GEN_95) : $signed(64'sh0); // @[Matrix_FixedPoint_Mul.scala 137:37 140:27 145:27]
  assign PE_FixedPoint_io_in_y = _T ? $signed(_GEN_211) : $signed(64'sh0); // @[Matrix_FixedPoint_Mul.scala 149:37 152:19 157:19]
  assign PE_FixedPoint_1_clock = clock;
  assign PE_FixedPoint_1_io_reset = io_reset | io_ready; // @[Matrix_FixedPoint_Mul.scala 85:18 95:20]
  assign PE_FixedPoint_1_io_in_x = PE_FixedPoint_io_out_x; // @[Matrix_FixedPoint_Mul.scala 167:17]
  assign PE_FixedPoint_1_io_in_y = _T ? $signed(_GEN_239) : $signed(64'sh0); // @[Matrix_FixedPoint_Mul.scala 149:37 152:19 157:19]
  assign PE_FixedPoint_2_clock = clock;
  assign PE_FixedPoint_2_io_reset = io_reset | io_ready; // @[Matrix_FixedPoint_Mul.scala 85:18 95:20]
  assign PE_FixedPoint_2_io_in_x = PE_FixedPoint_1_io_out_x; // @[Matrix_FixedPoint_Mul.scala 167:17]
  assign PE_FixedPoint_2_io_in_y = _T ? $signed(_GEN_267) : $signed(64'sh0); // @[Matrix_FixedPoint_Mul.scala 149:37 152:19 157:19]
  assign PE_FixedPoint_3_clock = clock;
  assign PE_FixedPoint_3_io_reset = io_reset | io_ready; // @[Matrix_FixedPoint_Mul.scala 85:18 95:20]
  assign PE_FixedPoint_3_io_in_x = PE_FixedPoint_2_io_out_x; // @[Matrix_FixedPoint_Mul.scala 167:17]
  assign PE_FixedPoint_3_io_in_y = _T ? $signed(_GEN_295) : $signed(64'sh0); // @[Matrix_FixedPoint_Mul.scala 149:37 152:19 157:19]
  assign PE_FixedPoint_4_clock = clock;
  assign PE_FixedPoint_4_io_reset = io_reset | io_ready; // @[Matrix_FixedPoint_Mul.scala 85:18 95:20]
  assign PE_FixedPoint_4_io_in_x = input_point < 5'h7 ? $signed(_GEN_123) : $signed(64'sh0); // @[Matrix_FixedPoint_Mul.scala 137:37 140:27 145:27]
  assign PE_FixedPoint_4_io_in_y = PE_FixedPoint_io_out_y; // @[Matrix_FixedPoint_Mul.scala 164:25]
  assign PE_FixedPoint_5_clock = clock;
  assign PE_FixedPoint_5_io_reset = io_reset | io_ready; // @[Matrix_FixedPoint_Mul.scala 85:18 95:20]
  assign PE_FixedPoint_5_io_in_x = PE_FixedPoint_4_io_out_x; // @[Matrix_FixedPoint_Mul.scala 172:27]
  assign PE_FixedPoint_5_io_in_y = PE_FixedPoint_1_io_out_y; // @[Matrix_FixedPoint_Mul.scala 171:27]
  assign PE_FixedPoint_6_clock = clock;
  assign PE_FixedPoint_6_io_reset = io_reset | io_ready; // @[Matrix_FixedPoint_Mul.scala 85:18 95:20]
  assign PE_FixedPoint_6_io_in_x = PE_FixedPoint_5_io_out_x; // @[Matrix_FixedPoint_Mul.scala 172:27]
  assign PE_FixedPoint_6_io_in_y = PE_FixedPoint_2_io_out_y; // @[Matrix_FixedPoint_Mul.scala 171:27]
  assign PE_FixedPoint_7_clock = clock;
  assign PE_FixedPoint_7_io_reset = io_reset | io_ready; // @[Matrix_FixedPoint_Mul.scala 85:18 95:20]
  assign PE_FixedPoint_7_io_in_x = PE_FixedPoint_6_io_out_x; // @[Matrix_FixedPoint_Mul.scala 172:27]
  assign PE_FixedPoint_7_io_in_y = PE_FixedPoint_3_io_out_y; // @[Matrix_FixedPoint_Mul.scala 171:27]
  assign PE_FixedPoint_8_clock = clock;
  assign PE_FixedPoint_8_io_reset = io_reset | io_ready; // @[Matrix_FixedPoint_Mul.scala 85:18 95:20]
  assign PE_FixedPoint_8_io_in_x = input_point < 5'h7 ? $signed(_GEN_151) : $signed(64'sh0); // @[Matrix_FixedPoint_Mul.scala 137:37 140:27 145:27]
  assign PE_FixedPoint_8_io_in_y = PE_FixedPoint_4_io_out_y; // @[Matrix_FixedPoint_Mul.scala 164:25]
  assign PE_FixedPoint_9_clock = clock;
  assign PE_FixedPoint_9_io_reset = io_reset | io_ready; // @[Matrix_FixedPoint_Mul.scala 85:18 95:20]
  assign PE_FixedPoint_9_io_in_x = PE_FixedPoint_8_io_out_x; // @[Matrix_FixedPoint_Mul.scala 172:27]
  assign PE_FixedPoint_9_io_in_y = PE_FixedPoint_5_io_out_y; // @[Matrix_FixedPoint_Mul.scala 171:27]
  assign PE_FixedPoint_10_clock = clock;
  assign PE_FixedPoint_10_io_reset = io_reset | io_ready; // @[Matrix_FixedPoint_Mul.scala 85:18 95:20]
  assign PE_FixedPoint_10_io_in_x = PE_FixedPoint_9_io_out_x; // @[Matrix_FixedPoint_Mul.scala 172:27]
  assign PE_FixedPoint_10_io_in_y = PE_FixedPoint_6_io_out_y; // @[Matrix_FixedPoint_Mul.scala 171:27]
  assign PE_FixedPoint_11_clock = clock;
  assign PE_FixedPoint_11_io_reset = io_reset | io_ready; // @[Matrix_FixedPoint_Mul.scala 85:18 95:20]
  assign PE_FixedPoint_11_io_in_x = PE_FixedPoint_10_io_out_x; // @[Matrix_FixedPoint_Mul.scala 172:27]
  assign PE_FixedPoint_11_io_in_y = PE_FixedPoint_7_io_out_y; // @[Matrix_FixedPoint_Mul.scala 171:27]
  assign PE_FixedPoint_12_clock = clock;
  assign PE_FixedPoint_12_io_reset = io_reset | io_ready; // @[Matrix_FixedPoint_Mul.scala 85:18 95:20]
  assign PE_FixedPoint_12_io_in_x = input_point < 5'h7 ? $signed(_GEN_179) : $signed(64'sh0); // @[Matrix_FixedPoint_Mul.scala 137:37 140:27 145:27]
  assign PE_FixedPoint_12_io_in_y = PE_FixedPoint_8_io_out_y; // @[Matrix_FixedPoint_Mul.scala 164:25]
  assign PE_FixedPoint_13_clock = clock;
  assign PE_FixedPoint_13_io_reset = io_reset | io_ready; // @[Matrix_FixedPoint_Mul.scala 85:18 95:20]
  assign PE_FixedPoint_13_io_in_x = PE_FixedPoint_12_io_out_x; // @[Matrix_FixedPoint_Mul.scala 172:27]
  assign PE_FixedPoint_13_io_in_y = PE_FixedPoint_9_io_out_y; // @[Matrix_FixedPoint_Mul.scala 171:27]
  assign PE_FixedPoint_14_clock = clock;
  assign PE_FixedPoint_14_io_reset = io_reset | io_ready; // @[Matrix_FixedPoint_Mul.scala 85:18 95:20]
  assign PE_FixedPoint_14_io_in_x = PE_FixedPoint_13_io_out_x; // @[Matrix_FixedPoint_Mul.scala 172:27]
  assign PE_FixedPoint_14_io_in_y = PE_FixedPoint_10_io_out_y; // @[Matrix_FixedPoint_Mul.scala 171:27]
  assign PE_FixedPoint_15_clock = clock;
  assign PE_FixedPoint_15_io_reset = io_reset | io_ready; // @[Matrix_FixedPoint_Mul.scala 85:18 95:20]
  assign PE_FixedPoint_15_io_in_x = PE_FixedPoint_14_io_out_x; // @[Matrix_FixedPoint_Mul.scala 172:27]
  assign PE_FixedPoint_15_io_in_y = PE_FixedPoint_11_io_out_y; // @[Matrix_FixedPoint_Mul.scala 171:27]
  always @(posedge clock) begin
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsA_0 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 88:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsA_0 <= io_matrixA_0; // @[Matrix_FixedPoint_Mul.scala 99:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsA_4 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 88:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsA_4 <= io_matrixA_4; // @[Matrix_FixedPoint_Mul.scala 99:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsA_5 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 88:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsA_5 <= io_matrixA_5; // @[Matrix_FixedPoint_Mul.scala 99:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsA_8 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 88:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsA_8 <= io_matrixA_8; // @[Matrix_FixedPoint_Mul.scala 99:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsA_9 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 88:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsA_9 <= io_matrixA_9; // @[Matrix_FixedPoint_Mul.scala 99:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsA_10 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 88:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsA_10 <= io_matrixA_10; // @[Matrix_FixedPoint_Mul.scala 99:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsA_12 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 88:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsA_12 <= io_matrixA_12; // @[Matrix_FixedPoint_Mul.scala 99:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsA_13 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 88:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsA_13 <= io_matrixA_13; // @[Matrix_FixedPoint_Mul.scala 99:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsA_14 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 88:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsA_14 <= io_matrixA_14; // @[Matrix_FixedPoint_Mul.scala 99:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsA_15 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 88:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsA_15 <= io_matrixA_15; // @[Matrix_FixedPoint_Mul.scala 99:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsB_0 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 91:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsB_0 <= io_matrixB_0; // @[Matrix_FixedPoint_Mul.scala 100:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsB_4 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 91:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsB_4 <= io_matrixB_4; // @[Matrix_FixedPoint_Mul.scala 100:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsB_5 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 91:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsB_5 <= io_matrixB_5; // @[Matrix_FixedPoint_Mul.scala 100:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsB_8 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 91:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsB_8 <= io_matrixB_8; // @[Matrix_FixedPoint_Mul.scala 100:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsB_9 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 91:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsB_9 <= io_matrixB_9; // @[Matrix_FixedPoint_Mul.scala 100:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsB_10 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 91:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsB_10 <= io_matrixB_10; // @[Matrix_FixedPoint_Mul.scala 100:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsB_12 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 91:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsB_12 <= io_matrixB_12; // @[Matrix_FixedPoint_Mul.scala 100:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsB_13 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 91:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsB_13 <= io_matrixB_13; // @[Matrix_FixedPoint_Mul.scala 100:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsB_14 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 91:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsB_14 <= io_matrixB_14; // @[Matrix_FixedPoint_Mul.scala 100:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      regsB_15 <= 64'sh0; // @[Matrix_FixedPoint_Mul.scala 91:16]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      regsB_15 <= io_matrixB_15; // @[Matrix_FixedPoint_Mul.scala 100:11]
    end
    if (io_reset) begin // @[Matrix_FixedPoint_Mul.scala 85:18]
      input_point <= 5'h0; // @[Matrix_FixedPoint_Mul.scala 93:17]
    end else if (io_ready) begin // @[Matrix_FixedPoint_Mul.scala 97:24]
      input_point <= 5'h0; // @[Matrix_FixedPoint_Mul.scala 102:17]
    end else begin
      input_point <= _input_point_T_1; // @[Matrix_FixedPoint_Mul.scala 110:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regsA_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regsA_4 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  regsA_5 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  regsA_8 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  regsA_9 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  regsA_10 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  regsA_12 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  regsA_13 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  regsA_14 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  regsA_15 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  regsB_0 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  regsB_4 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  regsB_5 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  regsB_8 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  regsB_9 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  regsB_10 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  regsB_12 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  regsB_13 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  regsB_14 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  regsB_15 = _RAND_19[63:0];
  _RAND_20 = {1{`RANDOM}};
  input_point = _RAND_20[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module mac_fixedpoint_v1(
  input  [63:0] io_vectorA_0,
  input  [63:0] io_vectorB_0,
  output [63:0] io_result
);
  wire [127:0] _res_0_T = $signed(io_vectorA_0) * $signed(io_vectorB_0); // @[Lower_Triangular_Matrix_Inversion_V1.scala 25:31]
  wire [95:0] _GEN_0 = _res_0_T[127:32]; // @[Lower_Triangular_Matrix_Inversion_V1.scala 21:17 25:14]
  assign io_result = _GEN_0[63:0]; // @[Lower_Triangular_Matrix_Inversion_V1.scala 21:17 25:14]
endmodule
module mac_fixedpoint_v1_3(
  input  [63:0] io_vectorA_0,
  input  [63:0] io_vectorA_1,
  input  [63:0] io_vectorB_0,
  input  [63:0] io_vectorB_1,
  output [63:0] io_result
);
  wire [127:0] _res_0_T = $signed(io_vectorA_0) * $signed(io_vectorB_0); // @[Lower_Triangular_Matrix_Inversion_V1.scala 25:31]
  wire [127:0] _res_1_T = $signed(io_vectorA_1) * $signed(io_vectorB_1); // @[Lower_Triangular_Matrix_Inversion_V1.scala 27:44]
  wire [95:0] _GEN_0 = _res_0_T[127:32]; // @[Lower_Triangular_Matrix_Inversion_V1.scala 21:17 25:14]
  wire [63:0] res_0 = _GEN_0[63:0]; // @[Lower_Triangular_Matrix_Inversion_V1.scala 21:17 25:14]
  wire [95:0] _GEN_2 = {$signed(res_0), 32'h0}; // @[Lower_Triangular_Matrix_Inversion_V1.scala 27:28]
  wire [127:0] _GEN_3 = {{32{_GEN_2[95]}},_GEN_2}; // @[Lower_Triangular_Matrix_Inversion_V1.scala 27:28]
  wire [127:0] _res_1_T_3 = $signed(_GEN_3) + $signed(_res_1_T); // @[Lower_Triangular_Matrix_Inversion_V1.scala 27:28]
  wire [95:0] _GEN_4 = _res_1_T_3[127:32]; // @[Lower_Triangular_Matrix_Inversion_V1.scala 21:17 27:14]
  assign io_result = _GEN_4[63:0]; // @[Lower_Triangular_Matrix_Inversion_V1.scala 21:17 27:14]
endmodule
module mac_fixedpoint_v1_5(
  input  [63:0] io_vectorA_0,
  input  [63:0] io_vectorA_1,
  input  [63:0] io_vectorA_2,
  input  [63:0] io_vectorB_0,
  input  [63:0] io_vectorB_1,
  input  [63:0] io_vectorB_2,
  output [63:0] io_result
);
  wire [127:0] _res_0_T = $signed(io_vectorA_0) * $signed(io_vectorB_0); // @[Lower_Triangular_Matrix_Inversion_V1.scala 25:31]
  wire [127:0] _res_1_T = $signed(io_vectorA_1) * $signed(io_vectorB_1); // @[Lower_Triangular_Matrix_Inversion_V1.scala 27:44]
  wire [95:0] _GEN_0 = _res_0_T[127:32]; // @[Lower_Triangular_Matrix_Inversion_V1.scala 21:17 25:14]
  wire [63:0] res_0 = _GEN_0[63:0]; // @[Lower_Triangular_Matrix_Inversion_V1.scala 21:17 25:14]
  wire [95:0] _GEN_2 = {$signed(res_0), 32'h0}; // @[Lower_Triangular_Matrix_Inversion_V1.scala 27:28]
  wire [127:0] _GEN_3 = {{32{_GEN_2[95]}},_GEN_2}; // @[Lower_Triangular_Matrix_Inversion_V1.scala 27:28]
  wire [127:0] _res_1_T_3 = $signed(_GEN_3) + $signed(_res_1_T); // @[Lower_Triangular_Matrix_Inversion_V1.scala 27:28]
  wire [127:0] _res_2_T = $signed(io_vectorA_2) * $signed(io_vectorB_2); // @[Lower_Triangular_Matrix_Inversion_V1.scala 27:44]
  wire [95:0] _GEN_4 = _res_1_T_3[127:32]; // @[Lower_Triangular_Matrix_Inversion_V1.scala 21:17 27:14]
  wire [63:0] res_1 = _GEN_4[63:0]; // @[Lower_Triangular_Matrix_Inversion_V1.scala 21:17 27:14]
  wire [95:0] _GEN_6 = {$signed(res_1), 32'h0}; // @[Lower_Triangular_Matrix_Inversion_V1.scala 27:28]
  wire [127:0] _GEN_7 = {{32{_GEN_6[95]}},_GEN_6}; // @[Lower_Triangular_Matrix_Inversion_V1.scala 27:28]
  wire [127:0] _res_2_T_3 = $signed(_GEN_7) + $signed(_res_2_T); // @[Lower_Triangular_Matrix_Inversion_V1.scala 27:28]
  wire [95:0] _GEN_8 = _res_2_T_3[127:32]; // @[Lower_Triangular_Matrix_Inversion_V1.scala 21:17 27:14]
  assign io_result = _GEN_8[63:0]; // @[Lower_Triangular_Matrix_Inversion_V1.scala 21:17 27:14]
endmodule
module lower_triangular_matrix_inversion_fixedpoint_v1(
  input         clock,
  input         reset,
  input         io_reset,
  input         io_ready,
  input  [63:0] io_matrixIn_0,
  input  [63:0] io_matrixIn_1,
  input  [63:0] io_matrixIn_2,
  input  [63:0] io_matrixIn_3,
  input  [63:0] io_matrixIn_4,
  input  [63:0] io_matrixIn_5,
  input  [63:0] io_matrixIn_6,
  input  [63:0] io_matrixIn_7,
  input  [63:0] io_matrixIn_8,
  input  [63:0] io_matrixIn_9,
  output [63:0] io_matrixOut_0,
  output [63:0] io_matrixOut_1,
  output [63:0] io_matrixOut_2,
  output [63:0] io_matrixOut_3,
  output [63:0] io_matrixOut_4,
  output [63:0] io_matrixOut_5,
  output [63:0] io_matrixOut_6,
  output [63:0] io_matrixOut_7,
  output [63:0] io_matrixOut_8,
  output [63:0] io_matrixOut_9,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire  reg_out_0_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  reg_out_0_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_0_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_0_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_0_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  reg_out_2_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  reg_out_2_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_2_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_2_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_2_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  reg_out_5_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  reg_out_5_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_5_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_5_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_5_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire  reg_out_9_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  reg_out_9_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_9_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_9_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_9_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire [63:0] mac_res_unit_io_vectorA_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_io_vectorB_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_io_result; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire  reg_out_1_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  reg_out_1_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_1_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_1_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_1_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire [63:0] mac_res_unit_1_io_vectorA_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_1_io_vectorB_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_1_io_result; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire  reg_out_4_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  reg_out_4_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_4_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_4_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_4_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire [63:0] mac_res_unit_2_io_vectorA_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_2_io_vectorB_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_2_io_result; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire  reg_out_8_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  reg_out_8_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_8_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_8_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_8_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire [63:0] mac_res_unit_3_io_vectorA_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_3_io_vectorA_1; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_3_io_vectorB_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_3_io_vectorB_1; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_3_io_result; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire  reg_out_3_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  reg_out_3_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_3_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_3_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_3_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire [63:0] mac_res_unit_4_io_vectorA_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_4_io_vectorA_1; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_4_io_vectorB_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_4_io_vectorB_1; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_4_io_result; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire  reg_out_7_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  reg_out_7_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_7_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_7_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_7_divide_io_z; // @[Cordic_LV.scala 211:24]
  wire [63:0] mac_res_unit_5_io_vectorA_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_5_io_vectorA_1; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_5_io_vectorA_2; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_5_io_vectorB_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_5_io_vectorB_1; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_5_io_vectorB_2; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire [63:0] mac_res_unit_5_io_result; // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
  wire  reg_out_6_divide_clock; // @[Cordic_LV.scala 211:24]
  wire  reg_out_6_divide_reset; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_6_divide_io_x; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_6_divide_io_y; // @[Cordic_LV.scala 211:24]
  wire [63:0] reg_out_6_divide_io_z; // @[Cordic_LV.scala 211:24]
  reg [63:0] reg_in_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 76:36]
  reg [63:0] reg_in_1; // @[Lower_Triangular_Matrix_Inversion_V1.scala 76:36]
  reg [63:0] reg_in_2; // @[Lower_Triangular_Matrix_Inversion_V1.scala 76:36]
  reg [63:0] reg_in_3; // @[Lower_Triangular_Matrix_Inversion_V1.scala 76:36]
  reg [63:0] reg_in_4; // @[Lower_Triangular_Matrix_Inversion_V1.scala 76:36]
  reg [63:0] reg_in_5; // @[Lower_Triangular_Matrix_Inversion_V1.scala 76:36]
  reg [63:0] reg_in_6; // @[Lower_Triangular_Matrix_Inversion_V1.scala 76:36]
  reg [63:0] reg_in_7; // @[Lower_Triangular_Matrix_Inversion_V1.scala 76:36]
  reg [63:0] reg_in_8; // @[Lower_Triangular_Matrix_Inversion_V1.scala 76:36]
  reg [63:0] reg_in_9; // @[Lower_Triangular_Matrix_Inversion_V1.scala 76:36]
  reg [63:0] reg_out_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 77:37]
  reg [63:0] reg_out_1; // @[Lower_Triangular_Matrix_Inversion_V1.scala 77:37]
  reg [63:0] reg_out_2; // @[Lower_Triangular_Matrix_Inversion_V1.scala 77:37]
  reg [63:0] reg_out_3; // @[Lower_Triangular_Matrix_Inversion_V1.scala 77:37]
  reg [63:0] reg_out_4; // @[Lower_Triangular_Matrix_Inversion_V1.scala 77:37]
  reg [63:0] reg_out_5; // @[Lower_Triangular_Matrix_Inversion_V1.scala 77:37]
  reg [63:0] reg_out_6; // @[Lower_Triangular_Matrix_Inversion_V1.scala 77:37]
  reg [63:0] reg_out_7; // @[Lower_Triangular_Matrix_Inversion_V1.scala 77:37]
  reg [63:0] reg_out_8; // @[Lower_Triangular_Matrix_Inversion_V1.scala 77:37]
  reg [63:0] reg_out_9; // @[Lower_Triangular_Matrix_Inversion_V1.scala 77:37]
  reg [31:0] reg_clk_cnt; // @[Lower_Triangular_Matrix_Inversion_V1.scala 78:34]
  wire [31:0] _reg_clk_cnt_T_1 = reg_clk_cnt + 32'h1; // @[Lower_Triangular_Matrix_Inversion_V1.scala 92:32]
  cordic_divide reg_out_0_divide ( // @[Cordic_LV.scala 211:24]
    .clock(reg_out_0_divide_clock),
    .reset(reg_out_0_divide_reset),
    .io_x(reg_out_0_divide_io_x),
    .io_y(reg_out_0_divide_io_y),
    .io_z(reg_out_0_divide_io_z)
  );
  cordic_divide reg_out_2_divide ( // @[Cordic_LV.scala 211:24]
    .clock(reg_out_2_divide_clock),
    .reset(reg_out_2_divide_reset),
    .io_x(reg_out_2_divide_io_x),
    .io_y(reg_out_2_divide_io_y),
    .io_z(reg_out_2_divide_io_z)
  );
  cordic_divide reg_out_5_divide ( // @[Cordic_LV.scala 211:24]
    .clock(reg_out_5_divide_clock),
    .reset(reg_out_5_divide_reset),
    .io_x(reg_out_5_divide_io_x),
    .io_y(reg_out_5_divide_io_y),
    .io_z(reg_out_5_divide_io_z)
  );
  cordic_divide reg_out_9_divide ( // @[Cordic_LV.scala 211:24]
    .clock(reg_out_9_divide_clock),
    .reset(reg_out_9_divide_reset),
    .io_x(reg_out_9_divide_io_x),
    .io_y(reg_out_9_divide_io_y),
    .io_z(reg_out_9_divide_io_z)
  );
  mac_fixedpoint_v1 mac_res_unit ( // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
    .io_vectorA_0(mac_res_unit_io_vectorA_0),
    .io_vectorB_0(mac_res_unit_io_vectorB_0),
    .io_result(mac_res_unit_io_result)
  );
  cordic_divide reg_out_1_divide ( // @[Cordic_LV.scala 211:24]
    .clock(reg_out_1_divide_clock),
    .reset(reg_out_1_divide_reset),
    .io_x(reg_out_1_divide_io_x),
    .io_y(reg_out_1_divide_io_y),
    .io_z(reg_out_1_divide_io_z)
  );
  mac_fixedpoint_v1 mac_res_unit_1 ( // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
    .io_vectorA_0(mac_res_unit_1_io_vectorA_0),
    .io_vectorB_0(mac_res_unit_1_io_vectorB_0),
    .io_result(mac_res_unit_1_io_result)
  );
  cordic_divide reg_out_4_divide ( // @[Cordic_LV.scala 211:24]
    .clock(reg_out_4_divide_clock),
    .reset(reg_out_4_divide_reset),
    .io_x(reg_out_4_divide_io_x),
    .io_y(reg_out_4_divide_io_y),
    .io_z(reg_out_4_divide_io_z)
  );
  mac_fixedpoint_v1 mac_res_unit_2 ( // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
    .io_vectorA_0(mac_res_unit_2_io_vectorA_0),
    .io_vectorB_0(mac_res_unit_2_io_vectorB_0),
    .io_result(mac_res_unit_2_io_result)
  );
  cordic_divide reg_out_8_divide ( // @[Cordic_LV.scala 211:24]
    .clock(reg_out_8_divide_clock),
    .reset(reg_out_8_divide_reset),
    .io_x(reg_out_8_divide_io_x),
    .io_y(reg_out_8_divide_io_y),
    .io_z(reg_out_8_divide_io_z)
  );
  mac_fixedpoint_v1_3 mac_res_unit_3 ( // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
    .io_vectorA_0(mac_res_unit_3_io_vectorA_0),
    .io_vectorA_1(mac_res_unit_3_io_vectorA_1),
    .io_vectorB_0(mac_res_unit_3_io_vectorB_0),
    .io_vectorB_1(mac_res_unit_3_io_vectorB_1),
    .io_result(mac_res_unit_3_io_result)
  );
  cordic_divide reg_out_3_divide ( // @[Cordic_LV.scala 211:24]
    .clock(reg_out_3_divide_clock),
    .reset(reg_out_3_divide_reset),
    .io_x(reg_out_3_divide_io_x),
    .io_y(reg_out_3_divide_io_y),
    .io_z(reg_out_3_divide_io_z)
  );
  mac_fixedpoint_v1_3 mac_res_unit_4 ( // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
    .io_vectorA_0(mac_res_unit_4_io_vectorA_0),
    .io_vectorA_1(mac_res_unit_4_io_vectorA_1),
    .io_vectorB_0(mac_res_unit_4_io_vectorB_0),
    .io_vectorB_1(mac_res_unit_4_io_vectorB_1),
    .io_result(mac_res_unit_4_io_result)
  );
  cordic_divide reg_out_7_divide ( // @[Cordic_LV.scala 211:24]
    .clock(reg_out_7_divide_clock),
    .reset(reg_out_7_divide_reset),
    .io_x(reg_out_7_divide_io_x),
    .io_y(reg_out_7_divide_io_y),
    .io_z(reg_out_7_divide_io_z)
  );
  mac_fixedpoint_v1_5 mac_res_unit_5 ( // @[Lower_Triangular_Matrix_Inversion_V1.scala 42:22]
    .io_vectorA_0(mac_res_unit_5_io_vectorA_0),
    .io_vectorA_1(mac_res_unit_5_io_vectorA_1),
    .io_vectorA_2(mac_res_unit_5_io_vectorA_2),
    .io_vectorB_0(mac_res_unit_5_io_vectorB_0),
    .io_vectorB_1(mac_res_unit_5_io_vectorB_1),
    .io_vectorB_2(mac_res_unit_5_io_vectorB_2),
    .io_result(mac_res_unit_5_io_result)
  );
  cordic_divide reg_out_6_divide ( // @[Cordic_LV.scala 211:24]
    .clock(reg_out_6_divide_clock),
    .reset(reg_out_6_divide_reset),
    .io_x(reg_out_6_divide_io_x),
    .io_y(reg_out_6_divide_io_y),
    .io_z(reg_out_6_divide_io_z)
  );
  assign io_matrixOut_0 = reg_out_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 130:16]
  assign io_matrixOut_1 = reg_out_1; // @[Lower_Triangular_Matrix_Inversion_V1.scala 130:16]
  assign io_matrixOut_2 = reg_out_2; // @[Lower_Triangular_Matrix_Inversion_V1.scala 130:16]
  assign io_matrixOut_3 = reg_out_3; // @[Lower_Triangular_Matrix_Inversion_V1.scala 130:16]
  assign io_matrixOut_4 = reg_out_4; // @[Lower_Triangular_Matrix_Inversion_V1.scala 130:16]
  assign io_matrixOut_5 = reg_out_5; // @[Lower_Triangular_Matrix_Inversion_V1.scala 130:16]
  assign io_matrixOut_6 = reg_out_6; // @[Lower_Triangular_Matrix_Inversion_V1.scala 130:16]
  assign io_matrixOut_7 = reg_out_7; // @[Lower_Triangular_Matrix_Inversion_V1.scala 130:16]
  assign io_matrixOut_8 = reg_out_8; // @[Lower_Triangular_Matrix_Inversion_V1.scala 130:16]
  assign io_matrixOut_9 = reg_out_9; // @[Lower_Triangular_Matrix_Inversion_V1.scala 130:16]
  assign io_valid = reg_clk_cnt >= 32'h40; // @[Lower_Triangular_Matrix_Inversion_V1.scala 125:20]
  assign reg_out_0_divide_clock = clock;
  assign reg_out_0_divide_reset = reset;
  assign reg_out_0_divide_io_x = reg_in_0; // @[Cordic_LV.scala 212:17]
  assign reg_out_0_divide_io_y = 64'sh100000000; // @[Cordic_LV.scala 213:17]
  assign reg_out_2_divide_clock = clock;
  assign reg_out_2_divide_reset = reset;
  assign reg_out_2_divide_io_x = reg_in_2; // @[Cordic_LV.scala 212:17]
  assign reg_out_2_divide_io_y = 64'sh100000000; // @[Cordic_LV.scala 213:17]
  assign reg_out_5_divide_clock = clock;
  assign reg_out_5_divide_reset = reset;
  assign reg_out_5_divide_io_x = reg_in_5; // @[Cordic_LV.scala 212:17]
  assign reg_out_5_divide_io_y = 64'sh100000000; // @[Cordic_LV.scala 213:17]
  assign reg_out_9_divide_clock = clock;
  assign reg_out_9_divide_reset = reset;
  assign reg_out_9_divide_io_x = reg_in_9; // @[Cordic_LV.scala 212:17]
  assign reg_out_9_divide_io_y = 64'sh100000000; // @[Cordic_LV.scala 213:17]
  assign mac_res_unit_io_vectorA_0 = reg_in_1; // @[Lower_Triangular_Matrix_Inversion_V1.scala 111:23 116:22]
  assign mac_res_unit_io_vectorB_0 = reg_out_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 112:23 117:22]
  assign reg_out_1_divide_clock = clock;
  assign reg_out_1_divide_reset = reset;
  assign reg_out_1_divide_io_x = reg_in_2; // @[Cordic_LV.scala 212:17]
  assign reg_out_1_divide_io_y = 64'sh0 - $signed(mac_res_unit_io_result); // @[Lower_Triangular_Matrix_Inversion_V1.scala 120:61]
  assign mac_res_unit_1_io_vectorA_0 = reg_in_4; // @[Lower_Triangular_Matrix_Inversion_V1.scala 111:23 116:22]
  assign mac_res_unit_1_io_vectorB_0 = reg_out_2; // @[Lower_Triangular_Matrix_Inversion_V1.scala 112:23 117:22]
  assign reg_out_4_divide_clock = clock;
  assign reg_out_4_divide_reset = reset;
  assign reg_out_4_divide_io_x = reg_in_5; // @[Cordic_LV.scala 212:17]
  assign reg_out_4_divide_io_y = 64'sh0 - $signed(mac_res_unit_1_io_result); // @[Lower_Triangular_Matrix_Inversion_V1.scala 120:61]
  assign mac_res_unit_2_io_vectorA_0 = reg_in_8; // @[Lower_Triangular_Matrix_Inversion_V1.scala 111:23 116:22]
  assign mac_res_unit_2_io_vectorB_0 = reg_out_5; // @[Lower_Triangular_Matrix_Inversion_V1.scala 112:23 117:22]
  assign reg_out_8_divide_clock = clock;
  assign reg_out_8_divide_reset = reset;
  assign reg_out_8_divide_io_x = reg_in_9; // @[Cordic_LV.scala 212:17]
  assign reg_out_8_divide_io_y = 64'sh0 - $signed(mac_res_unit_2_io_result); // @[Lower_Triangular_Matrix_Inversion_V1.scala 120:61]
  assign mac_res_unit_3_io_vectorA_0 = reg_in_3; // @[Lower_Triangular_Matrix_Inversion_V1.scala 111:23 116:22]
  assign mac_res_unit_3_io_vectorA_1 = reg_in_4; // @[Lower_Triangular_Matrix_Inversion_V1.scala 111:23 116:22]
  assign mac_res_unit_3_io_vectorB_0 = reg_out_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 112:23 117:22]
  assign mac_res_unit_3_io_vectorB_1 = reg_out_1; // @[Lower_Triangular_Matrix_Inversion_V1.scala 112:23 117:22]
  assign reg_out_3_divide_clock = clock;
  assign reg_out_3_divide_reset = reset;
  assign reg_out_3_divide_io_x = reg_in_5; // @[Cordic_LV.scala 212:17]
  assign reg_out_3_divide_io_y = 64'sh0 - $signed(mac_res_unit_3_io_result); // @[Lower_Triangular_Matrix_Inversion_V1.scala 120:61]
  assign mac_res_unit_4_io_vectorA_0 = reg_in_7; // @[Lower_Triangular_Matrix_Inversion_V1.scala 111:23 116:22]
  assign mac_res_unit_4_io_vectorA_1 = reg_in_8; // @[Lower_Triangular_Matrix_Inversion_V1.scala 111:23 116:22]
  assign mac_res_unit_4_io_vectorB_0 = reg_out_2; // @[Lower_Triangular_Matrix_Inversion_V1.scala 112:23 117:22]
  assign mac_res_unit_4_io_vectorB_1 = reg_out_4; // @[Lower_Triangular_Matrix_Inversion_V1.scala 112:23 117:22]
  assign reg_out_7_divide_clock = clock;
  assign reg_out_7_divide_reset = reset;
  assign reg_out_7_divide_io_x = reg_in_9; // @[Cordic_LV.scala 212:17]
  assign reg_out_7_divide_io_y = 64'sh0 - $signed(mac_res_unit_4_io_result); // @[Lower_Triangular_Matrix_Inversion_V1.scala 120:61]
  assign mac_res_unit_5_io_vectorA_0 = reg_in_6; // @[Lower_Triangular_Matrix_Inversion_V1.scala 111:23 116:22]
  assign mac_res_unit_5_io_vectorA_1 = reg_in_7; // @[Lower_Triangular_Matrix_Inversion_V1.scala 111:23 116:22]
  assign mac_res_unit_5_io_vectorA_2 = reg_in_8; // @[Lower_Triangular_Matrix_Inversion_V1.scala 111:23 116:22]
  assign mac_res_unit_5_io_vectorB_0 = reg_out_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 112:23 117:22]
  assign mac_res_unit_5_io_vectorB_1 = reg_out_1; // @[Lower_Triangular_Matrix_Inversion_V1.scala 112:23 117:22]
  assign mac_res_unit_5_io_vectorB_2 = reg_out_3; // @[Lower_Triangular_Matrix_Inversion_V1.scala 112:23 117:22]
  assign reg_out_6_divide_clock = clock;
  assign reg_out_6_divide_reset = reset;
  assign reg_out_6_divide_io_x = reg_in_9; // @[Cordic_LV.scala 212:17]
  assign reg_out_6_divide_io_y = 64'sh0 - $signed(mac_res_unit_5_io_result); // @[Lower_Triangular_Matrix_Inversion_V1.scala 120:61]
  always @(posedge clock) begin
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 81:18]
      reg_in_0 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 83:17]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 87:24]
      reg_in_0 <= io_matrixIn_0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 89:12]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 81:18]
      reg_in_1 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 83:17]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 87:24]
      reg_in_1 <= io_matrixIn_1; // @[Lower_Triangular_Matrix_Inversion_V1.scala 89:12]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 81:18]
      reg_in_2 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 83:17]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 87:24]
      reg_in_2 <= io_matrixIn_2; // @[Lower_Triangular_Matrix_Inversion_V1.scala 89:12]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 81:18]
      reg_in_3 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 83:17]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 87:24]
      reg_in_3 <= io_matrixIn_3; // @[Lower_Triangular_Matrix_Inversion_V1.scala 89:12]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 81:18]
      reg_in_4 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 83:17]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 87:24]
      reg_in_4 <= io_matrixIn_4; // @[Lower_Triangular_Matrix_Inversion_V1.scala 89:12]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 81:18]
      reg_in_5 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 83:17]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 87:24]
      reg_in_5 <= io_matrixIn_5; // @[Lower_Triangular_Matrix_Inversion_V1.scala 89:12]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 81:18]
      reg_in_6 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 83:17]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 87:24]
      reg_in_6 <= io_matrixIn_6; // @[Lower_Triangular_Matrix_Inversion_V1.scala 89:12]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 81:18]
      reg_in_7 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 83:17]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 87:24]
      reg_in_7 <= io_matrixIn_7; // @[Lower_Triangular_Matrix_Inversion_V1.scala 89:12]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 81:18]
      reg_in_8 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 83:17]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 87:24]
      reg_in_8 <= io_matrixIn_8; // @[Lower_Triangular_Matrix_Inversion_V1.scala 89:12]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 81:18]
      reg_in_9 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 83:17]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 87:24]
      reg_in_9 <= io_matrixIn_9; // @[Lower_Triangular_Matrix_Inversion_V1.scala 89:12]
    end
    reg_out_0 <= reg_out_0_divide_io_z; // @[Lower_Triangular_Matrix_Inversion_V1.scala 100:20]
    reg_out_1 <= reg_out_1_divide_io_z; // @[Lower_Triangular_Matrix_Inversion_V1.scala 120:26]
    reg_out_2 <= reg_out_2_divide_io_z; // @[Lower_Triangular_Matrix_Inversion_V1.scala 100:20]
    reg_out_3 <= reg_out_3_divide_io_z; // @[Lower_Triangular_Matrix_Inversion_V1.scala 120:26]
    reg_out_4 <= reg_out_4_divide_io_z; // @[Lower_Triangular_Matrix_Inversion_V1.scala 120:26]
    reg_out_5 <= reg_out_5_divide_io_z; // @[Lower_Triangular_Matrix_Inversion_V1.scala 100:20]
    reg_out_6 <= reg_out_6_divide_io_z; // @[Lower_Triangular_Matrix_Inversion_V1.scala 120:26]
    reg_out_7 <= reg_out_7_divide_io_z; // @[Lower_Triangular_Matrix_Inversion_V1.scala 120:26]
    reg_out_8 <= reg_out_8_divide_io_z; // @[Lower_Triangular_Matrix_Inversion_V1.scala 120:26]
    reg_out_9 <= reg_out_9_divide_io_z; // @[Lower_Triangular_Matrix_Inversion_V1.scala 100:20]
    if (reset) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 78:34]
      reg_clk_cnt <= 32'h0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 78:34]
    end else if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 81:18]
      reg_clk_cnt <= 32'h0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 86:17]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_V1.scala 87:24]
      reg_clk_cnt <= 32'h0; // @[Lower_Triangular_Matrix_Inversion_V1.scala 90:17]
    end else begin
      reg_clk_cnt <= _reg_clk_cnt_T_1; // @[Lower_Triangular_Matrix_Inversion_V1.scala 92:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  reg_in_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  reg_in_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  reg_in_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  reg_in_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  reg_in_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  reg_in_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  reg_in_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  reg_in_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  reg_in_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  reg_in_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  reg_out_0 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  reg_out_1 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  reg_out_2 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  reg_out_3 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  reg_out_4 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  reg_out_5 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  reg_out_6 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  reg_out_7 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  reg_out_8 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  reg_out_9 = _RAND_19[63:0];
  _RAND_20 = {1{`RANDOM}};
  reg_clk_cnt = _RAND_20[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module lower_triangular_matrix_inversion_complex_v1(
  input         clock,
  input         reset,
  input         io_reset,
  input         io_ready,
  input  [63:0] io_matrixIn_0_re,
  input  [63:0] io_matrixIn_0_im,
  input  [63:0] io_matrixIn_1_re,
  input  [63:0] io_matrixIn_1_im,
  input  [63:0] io_matrixIn_2_re,
  input  [63:0] io_matrixIn_2_im,
  input  [63:0] io_matrixIn_3_re,
  input  [63:0] io_matrixIn_3_im,
  input  [63:0] io_matrixIn_4_re,
  input  [63:0] io_matrixIn_4_im,
  input  [63:0] io_matrixIn_5_re,
  input  [63:0] io_matrixIn_5_im,
  input  [63:0] io_matrixIn_6_re,
  input  [63:0] io_matrixIn_6_im,
  input  [63:0] io_matrixIn_7_re,
  input  [63:0] io_matrixIn_7_im,
  input  [63:0] io_matrixIn_8_re,
  input  [63:0] io_matrixIn_8_im,
  input  [63:0] io_matrixIn_9_re,
  input  [63:0] io_matrixIn_9_im,
  output [63:0] io_matrixOut_0_re,
  output [63:0] io_matrixOut_0_im,
  output [63:0] io_matrixOut_1_re,
  output [63:0] io_matrixOut_1_im,
  output [63:0] io_matrixOut_2_re,
  output [63:0] io_matrixOut_2_im,
  output [63:0] io_matrixOut_3_re,
  output [63:0] io_matrixOut_3_im,
  output [63:0] io_matrixOut_4_re,
  output [63:0] io_matrixOut_4_im,
  output [63:0] io_matrixOut_5_re,
  output [63:0] io_matrixOut_5_im,
  output [63:0] io_matrixOut_6_re,
  output [63:0] io_matrixOut_6_im,
  output [63:0] io_matrixOut_7_re,
  output [63:0] io_matrixOut_7_im,
  output [63:0] io_matrixOut_8_re,
  output [63:0] io_matrixOut_8_im,
  output [63:0] io_matrixOut_9_re,
  output [63:0] io_matrixOut_9_im,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [31:0] _RAND_60;
`endif // RANDOMIZE_REG_INIT
  wire  matrix_mul_unit_clock; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire  matrix_mul_unit_io_reset; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire  matrix_mul_unit_io_ready; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixA_0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixA_4; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixA_5; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixA_8; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixA_9; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixA_10; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixA_12; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixA_13; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixA_14; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixA_15; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixB_0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixB_4; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixB_5; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixB_8; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixB_9; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixB_10; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixB_12; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixB_13; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixB_14; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixB_15; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixC_0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixC_4; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixC_5; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixC_8; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixC_9; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixC_10; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixC_12; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixC_13; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixC_14; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire [63:0] matrix_mul_unit_io_matrixC_15; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire  matrix_mul_unit_io_valid; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
  wire  lower_tri_mat_inv_unit_clock; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire  lower_tri_mat_inv_unit_reset; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire  lower_tri_mat_inv_unit_io_reset; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire  lower_tri_mat_inv_unit_io_ready; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixIn_0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixIn_1; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixIn_2; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixIn_3; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixIn_4; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixIn_5; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixIn_6; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixIn_7; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixIn_8; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixIn_9; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixOut_0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixOut_1; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixOut_2; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixOut_3; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixOut_4; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixOut_5; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixOut_6; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixOut_7; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixOut_8; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire [63:0] lower_tri_mat_inv_unit_io_matrixOut_9; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  wire  lower_tri_mat_inv_unit_io_valid; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
  reg [63:0] reg_x_0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 36:35]
  reg [63:0] reg_x_1; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 36:35]
  reg [63:0] reg_x_2; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 36:35]
  reg [63:0] reg_x_3; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 36:35]
  reg [63:0] reg_x_4; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 36:35]
  reg [63:0] reg_x_5; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 36:35]
  reg [63:0] reg_x_6; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 36:35]
  reg [63:0] reg_x_7; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 36:35]
  reg [63:0] reg_x_8; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 36:35]
  reg [63:0] reg_x_9; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 36:35]
  reg [63:0] reg_y_0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 37:35]
  reg [63:0] reg_y_1; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 37:35]
  reg [63:0] reg_y_2; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 37:35]
  reg [63:0] reg_y_3; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 37:35]
  reg [63:0] reg_y_4; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 37:35]
  reg [63:0] reg_y_5; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 37:35]
  reg [63:0] reg_y_6; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 37:35]
  reg [63:0] reg_y_7; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 37:35]
  reg [63:0] reg_y_8; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 37:35]
  reg [63:0] reg_y_9; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 37:35]
  reg [63:0] reg_x_inv_0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 38:39]
  reg [63:0] reg_x_inv_1; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 38:39]
  reg [63:0] reg_x_inv_2; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 38:39]
  reg [63:0] reg_x_inv_3; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 38:39]
  reg [63:0] reg_x_inv_4; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 38:39]
  reg [63:0] reg_x_inv_5; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 38:39]
  reg [63:0] reg_x_inv_6; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 38:39]
  reg [63:0] reg_x_inv_7; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 38:39]
  reg [63:0] reg_x_inv_8; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 38:39]
  reg [63:0] reg_x_inv_9; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 38:39]
  reg [63:0] reg_x_inv_y_0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 39:41]
  reg [63:0] reg_x_inv_y_1; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 39:41]
  reg [63:0] reg_x_inv_y_2; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 39:41]
  reg [63:0] reg_x_inv_y_3; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 39:41]
  reg [63:0] reg_x_inv_y_4; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 39:41]
  reg [63:0] reg_x_inv_y_5; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 39:41]
  reg [63:0] reg_x_inv_y_6; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 39:41]
  reg [63:0] reg_x_inv_y_7; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 39:41]
  reg [63:0] reg_x_inv_y_8; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 39:41]
  reg [63:0] reg_x_inv_y_9; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 39:41]
  reg [63:0] reg_u_0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 40:35]
  reg [63:0] reg_u_1; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 40:35]
  reg [63:0] reg_u_2; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 40:35]
  reg [63:0] reg_u_3; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 40:35]
  reg [63:0] reg_u_4; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 40:35]
  reg [63:0] reg_u_5; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 40:35]
  reg [63:0] reg_u_6; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 40:35]
  reg [63:0] reg_u_7; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 40:35]
  reg [63:0] reg_u_8; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 40:35]
  reg [63:0] reg_u_9; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 40:35]
  reg [63:0] reg_v_0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 41:35]
  reg [63:0] reg_v_1; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 41:35]
  reg [63:0] reg_v_2; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 41:35]
  reg [63:0] reg_v_3; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 41:35]
  reg [63:0] reg_v_4; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 41:35]
  reg [63:0] reg_v_5; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 41:35]
  reg [63:0] reg_v_6; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 41:35]
  reg [63:0] reg_v_7; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 41:35]
  reg [63:0] reg_v_8; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 41:35]
  reg [63:0] reg_v_9; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 41:35]
  reg [3:0] reg_step_status; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 42:38]
  wire [3:0] _GEN_20 = io_ready ? 4'h1 : reg_step_status; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24 83:21 42:38]
  wire [63:0] _GEN_23 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_0); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 71:20 38:39]
  wire [63:0] _GEN_24 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_y_0); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 72:22 39:41]
  wire [63:0] _GEN_25 = io_reset ? $signed(64'sh0) : $signed(reg_u_0); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 73:16 40:35]
  wire [63:0] _GEN_26 = io_reset ? $signed(64'sh0) : $signed(reg_v_0); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 74:16 41:35]
  wire [63:0] _GEN_29 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_1); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 71:20 38:39]
  wire [63:0] _GEN_30 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_y_1); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 72:22 39:41]
  wire [63:0] _GEN_31 = io_reset ? $signed(64'sh0) : $signed(reg_u_1); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 73:16 40:35]
  wire [63:0] _GEN_32 = io_reset ? $signed(64'sh0) : $signed(reg_v_1); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 74:16 41:35]
  wire [63:0] _GEN_35 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 71:20 38:39]
  wire [63:0] _GEN_36 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_y_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 72:22 39:41]
  wire [63:0] _GEN_37 = io_reset ? $signed(64'sh0) : $signed(reg_u_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 73:16 40:35]
  wire [63:0] _GEN_38 = io_reset ? $signed(64'sh0) : $signed(reg_v_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 74:16 41:35]
  wire [63:0] _GEN_41 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_3); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 71:20 38:39]
  wire [63:0] _GEN_42 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_y_3); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 72:22 39:41]
  wire [63:0] _GEN_43 = io_reset ? $signed(64'sh0) : $signed(reg_u_3); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 73:16 40:35]
  wire [63:0] _GEN_44 = io_reset ? $signed(64'sh0) : $signed(reg_v_3); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 74:16 41:35]
  wire [63:0] _GEN_47 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_4); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 71:20 38:39]
  wire [63:0] _GEN_48 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_y_4); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 72:22 39:41]
  wire [63:0] _GEN_49 = io_reset ? $signed(64'sh0) : $signed(reg_u_4); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 73:16 40:35]
  wire [63:0] _GEN_50 = io_reset ? $signed(64'sh0) : $signed(reg_v_4); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 74:16 41:35]
  wire [63:0] _GEN_53 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_5); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 71:20 38:39]
  wire [63:0] _GEN_54 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_y_5); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 72:22 39:41]
  wire [63:0] _GEN_55 = io_reset ? $signed(64'sh0) : $signed(reg_u_5); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 73:16 40:35]
  wire [63:0] _GEN_56 = io_reset ? $signed(64'sh0) : $signed(reg_v_5); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 74:16 41:35]
  wire [63:0] _GEN_59 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_6); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 71:20 38:39]
  wire [63:0] _GEN_60 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_y_6); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 72:22 39:41]
  wire [63:0] _GEN_61 = io_reset ? $signed(64'sh0) : $signed(reg_u_6); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 73:16 40:35]
  wire [63:0] _GEN_62 = io_reset ? $signed(64'sh0) : $signed(reg_v_6); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 74:16 41:35]
  wire [63:0] _GEN_65 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_7); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 71:20 38:39]
  wire [63:0] _GEN_66 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_y_7); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 72:22 39:41]
  wire [63:0] _GEN_67 = io_reset ? $signed(64'sh0) : $signed(reg_u_7); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 73:16 40:35]
  wire [63:0] _GEN_68 = io_reset ? $signed(64'sh0) : $signed(reg_v_7); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 74:16 41:35]
  wire [63:0] _GEN_71 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_8); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 71:20 38:39]
  wire [63:0] _GEN_72 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_y_8); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 72:22 39:41]
  wire [63:0] _GEN_73 = io_reset ? $signed(64'sh0) : $signed(reg_u_8); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 73:16 40:35]
  wire [63:0] _GEN_74 = io_reset ? $signed(64'sh0) : $signed(reg_v_8); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 74:16 41:35]
  wire [63:0] _GEN_77 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_9); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 71:20 38:39]
  wire [63:0] _GEN_78 = io_reset ? $signed(64'sh0) : $signed(reg_x_inv_y_9); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 72:22 39:41]
  wire [63:0] _GEN_79 = io_reset ? $signed(64'sh0) : $signed(reg_u_9); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 73:16 40:35]
  wire [63:0] _GEN_80 = io_reset ? $signed(64'sh0) : $signed(reg_v_9); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 74:16 41:35]
  wire [3:0] _GEN_81 = io_reset ? 4'h0 : _GEN_20; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18 76:21]
  wire [3:0] _reg_step_status_T_1 = reg_step_status + 4'h1; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 90:40]
  wire [3:0] _GEN_82 = lower_tri_mat_inv_unit_io_valid ? _reg_step_status_T_1 : _GEN_81; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 94:43 96:23]
  wire [3:0] _GEN_93 = matrix_mul_unit_io_valid ? _reg_step_status_T_1 : _GEN_81; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 116:36 117:23]
  wire [63:0] _GEN_94 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_0) : $signed(_GEN_24); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 116:36 120:44]
  wire [63:0] _GEN_95 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_4) : $signed(_GEN_30); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 116:36 120:44]
  wire [63:0] _GEN_96 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_5) : $signed(_GEN_36); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 116:36 120:44]
  wire [63:0] _GEN_97 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_8) : $signed(_GEN_42); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 116:36 120:44]
  wire [63:0] _GEN_98 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_9) : $signed(_GEN_48); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 116:36 120:44]
  wire [63:0] _GEN_99 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_10) : $signed(_GEN_54); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 116:36 120:44]
  wire [63:0] _GEN_100 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_12) : $signed(_GEN_60); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 116:36 120:44]
  wire [63:0] _GEN_101 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_13) : $signed(_GEN_66); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 116:36 120:44]
  wire [63:0] _GEN_102 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_14) : $signed(_GEN_72); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 116:36 120:44]
  wire [63:0] _GEN_103 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_15) : $signed(_GEN_78); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 116:36 120:44]
  wire [63:0] _GEN_105 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_0) : $signed(_GEN_25); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 141:36 145:38]
  wire [63:0] _GEN_106 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_4) : $signed(_GEN_31); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 141:36 145:38]
  wire [63:0] _GEN_107 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_5) : $signed(_GEN_37); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 141:36 145:38]
  wire [63:0] _GEN_108 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_8) : $signed(_GEN_43); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 141:36 145:38]
  wire [63:0] _GEN_109 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_9) : $signed(_GEN_49); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 141:36 145:38]
  wire [63:0] _GEN_110 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_10) : $signed(_GEN_55); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 141:36 145:38]
  wire [63:0] _GEN_111 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_12) : $signed(_GEN_61); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 141:36 145:38]
  wire [63:0] _GEN_112 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_13) : $signed(_GEN_67); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 141:36 145:38]
  wire [63:0] _GEN_113 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_14) : $signed(_GEN_73); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 141:36 145:38]
  wire [63:0] _GEN_114 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_15) : $signed(_GEN_79); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 141:36 145:38]
  wire  _T_6 = reg_step_status == 4'h7; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:30]
  wire [63:0] temp_add_0 = $signed(reg_x_0) + $signed(reg_u_0); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 153:31]
  wire [63:0] temp_add_1 = $signed(reg_x_1) + $signed(reg_u_1); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 153:31]
  wire [63:0] temp_add_2 = $signed(reg_x_2) + $signed(reg_u_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 153:31]
  wire [63:0] temp_add_3 = $signed(reg_x_3) + $signed(reg_u_3); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 153:31]
  wire [63:0] temp_add_4 = $signed(reg_x_4) + $signed(reg_u_4); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 153:31]
  wire [63:0] temp_add_5 = $signed(reg_x_5) + $signed(reg_u_5); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 153:31]
  wire [63:0] temp_add_6 = $signed(reg_x_6) + $signed(reg_u_6); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 153:31]
  wire [63:0] temp_add_7 = $signed(reg_x_7) + $signed(reg_u_7); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 153:31]
  wire [63:0] temp_add_8 = $signed(reg_x_8) + $signed(reg_u_8); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 153:31]
  wire [63:0] temp_add_9 = $signed(reg_x_9) + $signed(reg_u_9); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 153:31]
  wire [63:0] _GEN_116 = lower_tri_mat_inv_unit_io_valid ? $signed(lower_tri_mat_inv_unit_io_matrixOut_0) : $signed(
    _GEN_25); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 161:43 164:13]
  wire [63:0] _GEN_117 = lower_tri_mat_inv_unit_io_valid ? $signed(lower_tri_mat_inv_unit_io_matrixOut_1) : $signed(
    _GEN_31); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 161:43 164:13]
  wire [63:0] _GEN_118 = lower_tri_mat_inv_unit_io_valid ? $signed(lower_tri_mat_inv_unit_io_matrixOut_2) : $signed(
    _GEN_37); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 161:43 164:13]
  wire [63:0] _GEN_119 = lower_tri_mat_inv_unit_io_valid ? $signed(lower_tri_mat_inv_unit_io_matrixOut_3) : $signed(
    _GEN_43); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 161:43 164:13]
  wire [63:0] _GEN_120 = lower_tri_mat_inv_unit_io_valid ? $signed(lower_tri_mat_inv_unit_io_matrixOut_4) : $signed(
    _GEN_49); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 161:43 164:13]
  wire [63:0] _GEN_121 = lower_tri_mat_inv_unit_io_valid ? $signed(lower_tri_mat_inv_unit_io_matrixOut_5) : $signed(
    _GEN_55); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 161:43 164:13]
  wire [63:0] _GEN_122 = lower_tri_mat_inv_unit_io_valid ? $signed(lower_tri_mat_inv_unit_io_matrixOut_6) : $signed(
    _GEN_61); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 161:43 164:13]
  wire [63:0] _GEN_123 = lower_tri_mat_inv_unit_io_valid ? $signed(lower_tri_mat_inv_unit_io_matrixOut_7) : $signed(
    _GEN_67); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 161:43 164:13]
  wire [63:0] _GEN_124 = lower_tri_mat_inv_unit_io_valid ? $signed(lower_tri_mat_inv_unit_io_matrixOut_8) : $signed(
    _GEN_73); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 161:43 164:13]
  wire [63:0] _GEN_125 = lower_tri_mat_inv_unit_io_valid ? $signed(lower_tri_mat_inv_unit_io_matrixOut_9) : $signed(
    _GEN_79); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 161:43 164:13]
  wire  _T_8 = reg_step_status == 4'h9; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 166:30]
  wire [63:0] _temp_matirxA_0_T_2 = 64'sh0 - $signed(reg_x_inv_y_0); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 175:36]
  wire [63:0] _temp_matirxA_4_T_2 = 64'sh0 - $signed(reg_x_inv_y_1); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 175:36]
  wire [63:0] _temp_matirxA_5_T_2 = 64'sh0 - $signed(reg_x_inv_y_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 175:36]
  wire [63:0] _temp_matirxA_8_T_2 = 64'sh0 - $signed(reg_x_inv_y_3); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 175:36]
  wire [63:0] _temp_matirxA_9_T_2 = 64'sh0 - $signed(reg_x_inv_y_4); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 175:36]
  wire [63:0] _temp_matirxA_10_T_2 = 64'sh0 - $signed(reg_x_inv_y_5); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 175:36]
  wire [63:0] _temp_matirxA_12_T_2 = 64'sh0 - $signed(reg_x_inv_y_6); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 175:36]
  wire [63:0] _temp_matirxA_13_T_2 = 64'sh0 - $signed(reg_x_inv_y_7); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 175:36]
  wire [63:0] _temp_matirxA_14_T_2 = 64'sh0 - $signed(reg_x_inv_y_8); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 175:36]
  wire [63:0] _temp_matirxA_15_T_2 = 64'sh0 - $signed(reg_x_inv_y_9); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 175:36]
  wire [63:0] _GEN_126 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_0) : $signed(_GEN_26); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 183:36 186:38]
  wire [63:0] _GEN_127 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_4) : $signed(_GEN_32); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 183:36 186:38]
  wire [63:0] _GEN_128 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_5) : $signed(_GEN_38); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 183:36 186:38]
  wire [63:0] _GEN_129 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_8) : $signed(_GEN_44); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 183:36 186:38]
  wire [63:0] _GEN_130 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_9) : $signed(_GEN_50); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 183:36 186:38]
  wire [63:0] _GEN_131 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_10) : $signed(_GEN_56); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 183:36 186:38]
  wire [63:0] _GEN_132 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_12) : $signed(_GEN_62); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 183:36 186:38]
  wire [63:0] _GEN_133 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_13) : $signed(_GEN_68); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 183:36 186:38]
  wire [63:0] _GEN_134 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_14) : $signed(_GEN_74); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 183:36 186:38]
  wire [63:0] _GEN_135 = matrix_mul_unit_io_valid ? $signed(matrix_mul_unit_io_matrixC_15) : $signed(_GEN_80); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 183:36 186:38]
  wire [63:0] _GEN_138 = reg_step_status == 4'ha ? $signed(_GEN_126) : $signed(_GEN_26); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 180:40]
  wire [63:0] _GEN_139 = reg_step_status == 4'ha ? $signed(_GEN_127) : $signed(_GEN_32); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 180:40]
  wire [63:0] _GEN_140 = reg_step_status == 4'ha ? $signed(_GEN_128) : $signed(_GEN_38); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 180:40]
  wire [63:0] _GEN_141 = reg_step_status == 4'ha ? $signed(_GEN_129) : $signed(_GEN_44); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 180:40]
  wire [63:0] _GEN_142 = reg_step_status == 4'ha ? $signed(_GEN_130) : $signed(_GEN_50); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 180:40]
  wire [63:0] _GEN_143 = reg_step_status == 4'ha ? $signed(_GEN_131) : $signed(_GEN_56); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 180:40]
  wire [63:0] _GEN_144 = reg_step_status == 4'ha ? $signed(_GEN_132) : $signed(_GEN_62); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 180:40]
  wire [63:0] _GEN_145 = reg_step_status == 4'ha ? $signed(_GEN_133) : $signed(_GEN_68); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 180:40]
  wire [63:0] _GEN_146 = reg_step_status == 4'ha ? $signed(_GEN_134) : $signed(_GEN_74); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 180:40]
  wire [63:0] _GEN_147 = reg_step_status == 4'ha ? $signed(_GEN_135) : $signed(_GEN_80); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 180:40]
  wire [3:0] _GEN_148 = reg_step_status == 4'ha ? _GEN_93 : _GEN_81; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 180:40]
  wire [3:0] _GEN_171 = reg_step_status == 4'h9 ? _reg_step_status_T_1 : _GEN_148; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 166:39 179:21]
  wire [63:0] _GEN_172 = reg_step_status == 4'h9 ? $signed(_GEN_26) : $signed(_GEN_138); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 166:39]
  wire [63:0] _GEN_173 = reg_step_status == 4'h9 ? $signed(_GEN_32) : $signed(_GEN_139); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 166:39]
  wire [63:0] _GEN_174 = reg_step_status == 4'h9 ? $signed(_GEN_38) : $signed(_GEN_140); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 166:39]
  wire [63:0] _GEN_175 = reg_step_status == 4'h9 ? $signed(_GEN_44) : $signed(_GEN_141); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 166:39]
  wire [63:0] _GEN_176 = reg_step_status == 4'h9 ? $signed(_GEN_50) : $signed(_GEN_142); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 166:39]
  wire [63:0] _GEN_177 = reg_step_status == 4'h9 ? $signed(_GEN_56) : $signed(_GEN_143); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 166:39]
  wire [63:0] _GEN_178 = reg_step_status == 4'h9 ? $signed(_GEN_62) : $signed(_GEN_144); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 166:39]
  wire [63:0] _GEN_179 = reg_step_status == 4'h9 ? $signed(_GEN_68) : $signed(_GEN_145); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 166:39]
  wire [63:0] _GEN_180 = reg_step_status == 4'h9 ? $signed(_GEN_74) : $signed(_GEN_146); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 166:39]
  wire [63:0] _GEN_181 = reg_step_status == 4'h9 ? $signed(_GEN_80) : $signed(_GEN_147); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 166:39]
  wire [3:0] _GEN_183 = reg_step_status == 4'h8 ? _GEN_82 : _GEN_171; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_184 = reg_step_status == 4'h8 ? $signed(_GEN_116) : $signed(_GEN_25); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_185 = reg_step_status == 4'h8 ? $signed(_GEN_117) : $signed(_GEN_31); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_186 = reg_step_status == 4'h8 ? $signed(_GEN_118) : $signed(_GEN_37); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_187 = reg_step_status == 4'h8 ? $signed(_GEN_119) : $signed(_GEN_43); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_188 = reg_step_status == 4'h8 ? $signed(_GEN_120) : $signed(_GEN_49); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_189 = reg_step_status == 4'h8 ? $signed(_GEN_121) : $signed(_GEN_55); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_190 = reg_step_status == 4'h8 ? $signed(_GEN_122) : $signed(_GEN_61); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_191 = reg_step_status == 4'h8 ? $signed(_GEN_123) : $signed(_GEN_67); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_192 = reg_step_status == 4'h8 ? $signed(_GEN_124) : $signed(_GEN_73); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_193 = reg_step_status == 4'h8 ? $signed(_GEN_125) : $signed(_GEN_79); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_216 = reg_step_status == 4'h8 ? $signed(_GEN_26) : $signed(_GEN_172); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_217 = reg_step_status == 4'h8 ? $signed(_GEN_32) : $signed(_GEN_173); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_218 = reg_step_status == 4'h8 ? $signed(_GEN_38) : $signed(_GEN_174); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_219 = reg_step_status == 4'h8 ? $signed(_GEN_44) : $signed(_GEN_175); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_220 = reg_step_status == 4'h8 ? $signed(_GEN_50) : $signed(_GEN_176); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_221 = reg_step_status == 4'h8 ? $signed(_GEN_56) : $signed(_GEN_177); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_222 = reg_step_status == 4'h8 ? $signed(_GEN_62) : $signed(_GEN_178); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_223 = reg_step_status == 4'h8 ? $signed(_GEN_68) : $signed(_GEN_179); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_224 = reg_step_status == 4'h8 ? $signed(_GEN_74) : $signed(_GEN_180); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [63:0] _GEN_225 = reg_step_status == 4'h8 ? $signed(_GEN_80) : $signed(_GEN_181); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 158:39]
  wire [3:0] _GEN_237 = reg_step_status == 4'h7 ? _reg_step_status_T_1 : _GEN_183; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39 157:21]
  wire [63:0] _GEN_238 = reg_step_status == 4'h7 ? $signed(_GEN_25) : $signed(_GEN_184); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_239 = reg_step_status == 4'h7 ? $signed(_GEN_31) : $signed(_GEN_185); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_240 = reg_step_status == 4'h7 ? $signed(_GEN_37) : $signed(_GEN_186); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_241 = reg_step_status == 4'h7 ? $signed(_GEN_43) : $signed(_GEN_187); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_242 = reg_step_status == 4'h7 ? $signed(_GEN_49) : $signed(_GEN_188); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_243 = reg_step_status == 4'h7 ? $signed(_GEN_55) : $signed(_GEN_189); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_244 = reg_step_status == 4'h7 ? $signed(_GEN_61) : $signed(_GEN_190); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_245 = reg_step_status == 4'h7 ? $signed(_GEN_67) : $signed(_GEN_191); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_246 = reg_step_status == 4'h7 ? $signed(_GEN_73) : $signed(_GEN_192); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_247 = reg_step_status == 4'h7 ? $signed(_GEN_79) : $signed(_GEN_193); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_270 = reg_step_status == 4'h7 ? $signed(_GEN_26) : $signed(_GEN_216); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_271 = reg_step_status == 4'h7 ? $signed(_GEN_32) : $signed(_GEN_217); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_272 = reg_step_status == 4'h7 ? $signed(_GEN_38) : $signed(_GEN_218); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_273 = reg_step_status == 4'h7 ? $signed(_GEN_44) : $signed(_GEN_219); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_274 = reg_step_status == 4'h7 ? $signed(_GEN_50) : $signed(_GEN_220); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_275 = reg_step_status == 4'h7 ? $signed(_GEN_56) : $signed(_GEN_221); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_276 = reg_step_status == 4'h7 ? $signed(_GEN_62) : $signed(_GEN_222); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_277 = reg_step_status == 4'h7 ? $signed(_GEN_68) : $signed(_GEN_223); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_278 = reg_step_status == 4'h7 ? $signed(_GEN_74) : $signed(_GEN_224); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire [63:0] _GEN_279 = reg_step_status == 4'h7 ? $signed(_GEN_80) : $signed(_GEN_225); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 149:39]
  wire  _GEN_280 = reg_step_status == 4'h6 ? 1'h0 : _T_8; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39 140:30]
  wire [3:0] _GEN_281 = reg_step_status == 4'h6 ? _GEN_93 : _GEN_237; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_282 = reg_step_status == 4'h6 ? $signed(_GEN_105) : $signed(_GEN_238); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_283 = reg_step_status == 4'h6 ? $signed(_GEN_106) : $signed(_GEN_239); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_284 = reg_step_status == 4'h6 ? $signed(_GEN_107) : $signed(_GEN_240); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_285 = reg_step_status == 4'h6 ? $signed(_GEN_108) : $signed(_GEN_241); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_286 = reg_step_status == 4'h6 ? $signed(_GEN_109) : $signed(_GEN_242); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_287 = reg_step_status == 4'h6 ? $signed(_GEN_110) : $signed(_GEN_243); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_288 = reg_step_status == 4'h6 ? $signed(_GEN_111) : $signed(_GEN_244); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_289 = reg_step_status == 4'h6 ? $signed(_GEN_112) : $signed(_GEN_245); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_290 = reg_step_status == 4'h6 ? $signed(_GEN_113) : $signed(_GEN_246); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_291 = reg_step_status == 4'h6 ? $signed(_GEN_114) : $signed(_GEN_247); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_324 = reg_step_status == 4'h6 ? $signed(_GEN_26) : $signed(_GEN_270); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_325 = reg_step_status == 4'h6 ? $signed(_GEN_32) : $signed(_GEN_271); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_326 = reg_step_status == 4'h6 ? $signed(_GEN_38) : $signed(_GEN_272); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_327 = reg_step_status == 4'h6 ? $signed(_GEN_44) : $signed(_GEN_273); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_328 = reg_step_status == 4'h6 ? $signed(_GEN_50) : $signed(_GEN_274); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_329 = reg_step_status == 4'h6 ? $signed(_GEN_56) : $signed(_GEN_275); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_330 = reg_step_status == 4'h6 ? $signed(_GEN_62) : $signed(_GEN_276); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_331 = reg_step_status == 4'h6 ? $signed(_GEN_68) : $signed(_GEN_277); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_332 = reg_step_status == 4'h6 ? $signed(_GEN_74) : $signed(_GEN_278); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire [63:0] _GEN_333 = reg_step_status == 4'h6 ? $signed(_GEN_80) : $signed(_GEN_279); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 138:39]
  wire  _GEN_334 = reg_step_status == 4'h5 | _GEN_280; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 126:30]
  wire [63:0] _GEN_335 = reg_step_status == 4'h5 ? $signed(reg_y_0) : $signed(_temp_matirxA_0_T_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 133:33]
  wire [63:0] _GEN_336 = reg_step_status == 4'h5 ? $signed(reg_x_inv_y_0) : $signed(reg_u_0); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 134:33]
  wire [63:0] _GEN_338 = reg_step_status == 4'h5 ? $signed(reg_y_1) : $signed(_temp_matirxA_4_T_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 133:33]
  wire [63:0] _GEN_339 = reg_step_status == 4'h5 ? $signed(reg_x_inv_y_1) : $signed(reg_u_1); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 134:33]
  wire [63:0] _GEN_340 = reg_step_status == 4'h5 ? $signed(reg_y_2) : $signed(_temp_matirxA_5_T_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 133:33]
  wire [63:0] _GEN_341 = reg_step_status == 4'h5 ? $signed(reg_x_inv_y_2) : $signed(reg_u_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 134:33]
  wire [63:0] _GEN_342 = reg_step_status == 4'h5 ? $signed(reg_y_3) : $signed(_temp_matirxA_8_T_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 133:33]
  wire [63:0] _GEN_343 = reg_step_status == 4'h5 ? $signed(reg_x_inv_y_3) : $signed(reg_u_3); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 134:33]
  wire [63:0] _GEN_344 = reg_step_status == 4'h5 ? $signed(reg_y_4) : $signed(_temp_matirxA_9_T_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 133:33]
  wire [63:0] _GEN_345 = reg_step_status == 4'h5 ? $signed(reg_x_inv_y_4) : $signed(reg_u_4); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 134:33]
  wire [63:0] _GEN_346 = reg_step_status == 4'h5 ? $signed(reg_y_5) : $signed(_temp_matirxA_10_T_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 133:33]
  wire [63:0] _GEN_347 = reg_step_status == 4'h5 ? $signed(reg_x_inv_y_5) : $signed(reg_u_5); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 134:33]
  wire [63:0] _GEN_348 = reg_step_status == 4'h5 ? $signed(reg_y_6) : $signed(_temp_matirxA_12_T_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 133:33]
  wire [63:0] _GEN_349 = reg_step_status == 4'h5 ? $signed(reg_x_inv_y_6) : $signed(reg_u_6); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 134:33]
  wire [63:0] _GEN_350 = reg_step_status == 4'h5 ? $signed(reg_y_7) : $signed(_temp_matirxA_13_T_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 133:33]
  wire [63:0] _GEN_351 = reg_step_status == 4'h5 ? $signed(reg_x_inv_y_7) : $signed(reg_u_7); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 134:33]
  wire [63:0] _GEN_352 = reg_step_status == 4'h5 ? $signed(reg_y_8) : $signed(_temp_matirxA_14_T_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 133:33]
  wire [63:0] _GEN_353 = reg_step_status == 4'h5 ? $signed(reg_x_inv_y_8) : $signed(reg_u_8); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 134:33]
  wire [63:0] _GEN_354 = reg_step_status == 4'h5 ? $signed(reg_y_9) : $signed(_temp_matirxA_15_T_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 133:33]
  wire [63:0] _GEN_355 = reg_step_status == 4'h5 ? $signed(reg_x_inv_y_9) : $signed(reg_u_9); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 134:33]
  wire [3:0] _GEN_356 = reg_step_status == 4'h5 ? _reg_step_status_T_1 : _GEN_281; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39 137:21]
  wire [63:0] _GEN_357 = reg_step_status == 4'h5 ? $signed(_GEN_25) : $signed(_GEN_282); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_358 = reg_step_status == 4'h5 ? $signed(_GEN_31) : $signed(_GEN_283); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_359 = reg_step_status == 4'h5 ? $signed(_GEN_37) : $signed(_GEN_284); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_360 = reg_step_status == 4'h5 ? $signed(_GEN_43) : $signed(_GEN_285); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_361 = reg_step_status == 4'h5 ? $signed(_GEN_49) : $signed(_GEN_286); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_362 = reg_step_status == 4'h5 ? $signed(_GEN_55) : $signed(_GEN_287); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_363 = reg_step_status == 4'h5 ? $signed(_GEN_61) : $signed(_GEN_288); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_364 = reg_step_status == 4'h5 ? $signed(_GEN_67) : $signed(_GEN_289); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_365 = reg_step_status == 4'h5 ? $signed(_GEN_73) : $signed(_GEN_290); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_366 = reg_step_status == 4'h5 ? $signed(_GEN_79) : $signed(_GEN_291); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_378 = reg_step_status == 4'h5 ? $signed(_GEN_26) : $signed(_GEN_324); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_379 = reg_step_status == 4'h5 ? $signed(_GEN_32) : $signed(_GEN_325); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_380 = reg_step_status == 4'h5 ? $signed(_GEN_38) : $signed(_GEN_326); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_381 = reg_step_status == 4'h5 ? $signed(_GEN_44) : $signed(_GEN_327); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_382 = reg_step_status == 4'h5 ? $signed(_GEN_50) : $signed(_GEN_328); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_383 = reg_step_status == 4'h5 ? $signed(_GEN_56) : $signed(_GEN_329); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_384 = reg_step_status == 4'h5 ? $signed(_GEN_62) : $signed(_GEN_330); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_385 = reg_step_status == 4'h5 ? $signed(_GEN_68) : $signed(_GEN_331); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_386 = reg_step_status == 4'h5 ? $signed(_GEN_74) : $signed(_GEN_332); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire [63:0] _GEN_387 = reg_step_status == 4'h5 ? $signed(_GEN_80) : $signed(_GEN_333); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 124:39]
  wire  _GEN_388 = reg_step_status == 4'h4 ? 1'h0 : _GEN_334; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39 115:30]
  wire [3:0] _GEN_389 = reg_step_status == 4'h4 ? _GEN_93 : _GEN_356; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
  wire  _GEN_516 = reg_step_status == 4'h2 ? 1'h0 : _T_6; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39 93:37]
  matrix_fixedPoint_mul matrix_mul_unit ( // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 44:31]
    .clock(matrix_mul_unit_clock),
    .io_reset(matrix_mul_unit_io_reset),
    .io_ready(matrix_mul_unit_io_ready),
    .io_matrixA_0(matrix_mul_unit_io_matrixA_0),
    .io_matrixA_4(matrix_mul_unit_io_matrixA_4),
    .io_matrixA_5(matrix_mul_unit_io_matrixA_5),
    .io_matrixA_8(matrix_mul_unit_io_matrixA_8),
    .io_matrixA_9(matrix_mul_unit_io_matrixA_9),
    .io_matrixA_10(matrix_mul_unit_io_matrixA_10),
    .io_matrixA_12(matrix_mul_unit_io_matrixA_12),
    .io_matrixA_13(matrix_mul_unit_io_matrixA_13),
    .io_matrixA_14(matrix_mul_unit_io_matrixA_14),
    .io_matrixA_15(matrix_mul_unit_io_matrixA_15),
    .io_matrixB_0(matrix_mul_unit_io_matrixB_0),
    .io_matrixB_4(matrix_mul_unit_io_matrixB_4),
    .io_matrixB_5(matrix_mul_unit_io_matrixB_5),
    .io_matrixB_8(matrix_mul_unit_io_matrixB_8),
    .io_matrixB_9(matrix_mul_unit_io_matrixB_9),
    .io_matrixB_10(matrix_mul_unit_io_matrixB_10),
    .io_matrixB_12(matrix_mul_unit_io_matrixB_12),
    .io_matrixB_13(matrix_mul_unit_io_matrixB_13),
    .io_matrixB_14(matrix_mul_unit_io_matrixB_14),
    .io_matrixB_15(matrix_mul_unit_io_matrixB_15),
    .io_matrixC_0(matrix_mul_unit_io_matrixC_0),
    .io_matrixC_4(matrix_mul_unit_io_matrixC_4),
    .io_matrixC_5(matrix_mul_unit_io_matrixC_5),
    .io_matrixC_8(matrix_mul_unit_io_matrixC_8),
    .io_matrixC_9(matrix_mul_unit_io_matrixC_9),
    .io_matrixC_10(matrix_mul_unit_io_matrixC_10),
    .io_matrixC_12(matrix_mul_unit_io_matrixC_12),
    .io_matrixC_13(matrix_mul_unit_io_matrixC_13),
    .io_matrixC_14(matrix_mul_unit_io_matrixC_14),
    .io_matrixC_15(matrix_mul_unit_io_matrixC_15),
    .io_valid(matrix_mul_unit_io_valid)
  );
  lower_triangular_matrix_inversion_fixedpoint_v1 lower_tri_mat_inv_unit ( // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 45:38]
    .clock(lower_tri_mat_inv_unit_clock),
    .reset(lower_tri_mat_inv_unit_reset),
    .io_reset(lower_tri_mat_inv_unit_io_reset),
    .io_ready(lower_tri_mat_inv_unit_io_ready),
    .io_matrixIn_0(lower_tri_mat_inv_unit_io_matrixIn_0),
    .io_matrixIn_1(lower_tri_mat_inv_unit_io_matrixIn_1),
    .io_matrixIn_2(lower_tri_mat_inv_unit_io_matrixIn_2),
    .io_matrixIn_3(lower_tri_mat_inv_unit_io_matrixIn_3),
    .io_matrixIn_4(lower_tri_mat_inv_unit_io_matrixIn_4),
    .io_matrixIn_5(lower_tri_mat_inv_unit_io_matrixIn_5),
    .io_matrixIn_6(lower_tri_mat_inv_unit_io_matrixIn_6),
    .io_matrixIn_7(lower_tri_mat_inv_unit_io_matrixIn_7),
    .io_matrixIn_8(lower_tri_mat_inv_unit_io_matrixIn_8),
    .io_matrixIn_9(lower_tri_mat_inv_unit_io_matrixIn_9),
    .io_matrixOut_0(lower_tri_mat_inv_unit_io_matrixOut_0),
    .io_matrixOut_1(lower_tri_mat_inv_unit_io_matrixOut_1),
    .io_matrixOut_2(lower_tri_mat_inv_unit_io_matrixOut_2),
    .io_matrixOut_3(lower_tri_mat_inv_unit_io_matrixOut_3),
    .io_matrixOut_4(lower_tri_mat_inv_unit_io_matrixOut_4),
    .io_matrixOut_5(lower_tri_mat_inv_unit_io_matrixOut_5),
    .io_matrixOut_6(lower_tri_mat_inv_unit_io_matrixOut_6),
    .io_matrixOut_7(lower_tri_mat_inv_unit_io_matrixOut_7),
    .io_matrixOut_8(lower_tri_mat_inv_unit_io_matrixOut_8),
    .io_matrixOut_9(lower_tri_mat_inv_unit_io_matrixOut_9),
    .io_valid(lower_tri_mat_inv_unit_io_valid)
  );
  assign io_matrixOut_0_re = reg_u_0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 200:24]
  assign io_matrixOut_0_im = reg_v_0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 201:24]
  assign io_matrixOut_1_re = reg_u_1; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 200:24]
  assign io_matrixOut_1_im = reg_v_1; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 201:24]
  assign io_matrixOut_2_re = reg_u_2; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 200:24]
  assign io_matrixOut_2_im = reg_v_2; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 201:24]
  assign io_matrixOut_3_re = reg_u_3; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 200:24]
  assign io_matrixOut_3_im = reg_v_3; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 201:24]
  assign io_matrixOut_4_re = reg_u_4; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 200:24]
  assign io_matrixOut_4_im = reg_v_4; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 201:24]
  assign io_matrixOut_5_re = reg_u_5; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 200:24]
  assign io_matrixOut_5_im = reg_v_5; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 201:24]
  assign io_matrixOut_6_re = reg_u_6; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 200:24]
  assign io_matrixOut_6_im = reg_v_6; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 201:24]
  assign io_matrixOut_7_re = reg_u_7; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 200:24]
  assign io_matrixOut_7_im = reg_v_7; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 201:24]
  assign io_matrixOut_8_re = reg_u_8; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 200:24]
  assign io_matrixOut_8_im = reg_v_8; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 201:24]
  assign io_matrixOut_9_re = reg_u_9; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 200:24]
  assign io_matrixOut_9_im = reg_v_9; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 201:24]
  assign io_valid = reg_step_status == 4'hb; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 193:24]
  assign matrix_mul_unit_clock = clock;
  assign matrix_mul_unit_io_reset = io_reset; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 46:28]
  assign matrix_mul_unit_io_ready = reg_step_status == 4'h3 | _GEN_388; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 101:30 99:39]
  assign matrix_mul_unit_io_matrixA_0 = reg_step_status == 4'h3 ? $signed(reg_x_inv_0) : $signed(_GEN_335); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 108:33 99:39]
  assign matrix_mul_unit_io_matrixA_4 = reg_step_status == 4'h3 ? $signed(reg_x_inv_1) : $signed(_GEN_338); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 108:33 99:39]
  assign matrix_mul_unit_io_matrixA_5 = reg_step_status == 4'h3 ? $signed(reg_x_inv_2) : $signed(_GEN_340); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 108:33 99:39]
  assign matrix_mul_unit_io_matrixA_8 = reg_step_status == 4'h3 ? $signed(reg_x_inv_3) : $signed(_GEN_342); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 108:33 99:39]
  assign matrix_mul_unit_io_matrixA_9 = reg_step_status == 4'h3 ? $signed(reg_x_inv_4) : $signed(_GEN_344); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 108:33 99:39]
  assign matrix_mul_unit_io_matrixA_10 = reg_step_status == 4'h3 ? $signed(reg_x_inv_5) : $signed(_GEN_346); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 108:33 99:39]
  assign matrix_mul_unit_io_matrixA_12 = reg_step_status == 4'h3 ? $signed(reg_x_inv_6) : $signed(_GEN_348); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 108:33 99:39]
  assign matrix_mul_unit_io_matrixA_13 = reg_step_status == 4'h3 ? $signed(reg_x_inv_7) : $signed(_GEN_350); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 108:33 99:39]
  assign matrix_mul_unit_io_matrixA_14 = reg_step_status == 4'h3 ? $signed(reg_x_inv_8) : $signed(_GEN_352); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 108:33 99:39]
  assign matrix_mul_unit_io_matrixA_15 = reg_step_status == 4'h3 ? $signed(reg_x_inv_9) : $signed(_GEN_354); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 108:33 99:39]
  assign matrix_mul_unit_io_matrixB_0 = reg_step_status == 4'h3 ? $signed(reg_y_0) : $signed(_GEN_336); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 109:33 99:39]
  assign matrix_mul_unit_io_matrixB_4 = reg_step_status == 4'h3 ? $signed(reg_y_1) : $signed(_GEN_339); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 109:33 99:39]
  assign matrix_mul_unit_io_matrixB_5 = reg_step_status == 4'h3 ? $signed(reg_y_2) : $signed(_GEN_341); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 109:33 99:39]
  assign matrix_mul_unit_io_matrixB_8 = reg_step_status == 4'h3 ? $signed(reg_y_3) : $signed(_GEN_343); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 109:33 99:39]
  assign matrix_mul_unit_io_matrixB_9 = reg_step_status == 4'h3 ? $signed(reg_y_4) : $signed(_GEN_345); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 109:33 99:39]
  assign matrix_mul_unit_io_matrixB_10 = reg_step_status == 4'h3 ? $signed(reg_y_5) : $signed(_GEN_347); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 109:33 99:39]
  assign matrix_mul_unit_io_matrixB_12 = reg_step_status == 4'h3 ? $signed(reg_y_6) : $signed(_GEN_349); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 109:33 99:39]
  assign matrix_mul_unit_io_matrixB_13 = reg_step_status == 4'h3 ? $signed(reg_y_7) : $signed(_GEN_351); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 109:33 99:39]
  assign matrix_mul_unit_io_matrixB_14 = reg_step_status == 4'h3 ? $signed(reg_y_8) : $signed(_GEN_353); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 109:33 99:39]
  assign matrix_mul_unit_io_matrixB_15 = reg_step_status == 4'h3 ? $signed(reg_y_9) : $signed(_GEN_355); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 109:33 99:39]
  assign lower_tri_mat_inv_unit_clock = clock;
  assign lower_tri_mat_inv_unit_reset = reset;
  assign lower_tri_mat_inv_unit_io_reset = io_reset; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 47:35]
  assign lower_tri_mat_inv_unit_io_ready = reg_step_status == 4'h1 | _GEN_516; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33 88:37]
  assign lower_tri_mat_inv_unit_io_matrixIn_0 = reg_step_status == 4'h1 ? $signed(reg_x_0) : $signed(temp_add_0); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33 89:40]
  assign lower_tri_mat_inv_unit_io_matrixIn_1 = reg_step_status == 4'h1 ? $signed(reg_x_1) : $signed(temp_add_1); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33 89:40]
  assign lower_tri_mat_inv_unit_io_matrixIn_2 = reg_step_status == 4'h1 ? $signed(reg_x_2) : $signed(temp_add_2); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33 89:40]
  assign lower_tri_mat_inv_unit_io_matrixIn_3 = reg_step_status == 4'h1 ? $signed(reg_x_3) : $signed(temp_add_3); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33 89:40]
  assign lower_tri_mat_inv_unit_io_matrixIn_4 = reg_step_status == 4'h1 ? $signed(reg_x_4) : $signed(temp_add_4); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33 89:40]
  assign lower_tri_mat_inv_unit_io_matrixIn_5 = reg_step_status == 4'h1 ? $signed(reg_x_5) : $signed(temp_add_5); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33 89:40]
  assign lower_tri_mat_inv_unit_io_matrixIn_6 = reg_step_status == 4'h1 ? $signed(reg_x_6) : $signed(temp_add_6); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33 89:40]
  assign lower_tri_mat_inv_unit_io_matrixIn_7 = reg_step_status == 4'h1 ? $signed(reg_x_7) : $signed(temp_add_7); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33 89:40]
  assign lower_tri_mat_inv_unit_io_matrixIn_8 = reg_step_status == 4'h1 ? $signed(reg_x_8) : $signed(temp_add_8); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33 89:40]
  assign lower_tri_mat_inv_unit_io_matrixIn_9 = reg_step_status == 4'h1 ? $signed(reg_x_9) : $signed(temp_add_9); // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33 89:40]
  always @(posedge clock) begin
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_x_0 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 69:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_x_0 <= io_matrixIn_0_re; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 80:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_x_1 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 69:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_x_1 <= io_matrixIn_1_re; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 80:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_x_2 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 69:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_x_2 <= io_matrixIn_2_re; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 80:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_x_3 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 69:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_x_3 <= io_matrixIn_3_re; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 80:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_x_4 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 69:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_x_4 <= io_matrixIn_4_re; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 80:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_x_5 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 69:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_x_5 <= io_matrixIn_5_re; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 80:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_x_6 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 69:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_x_6 <= io_matrixIn_6_re; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 80:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_x_7 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 69:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_x_7 <= io_matrixIn_7_re; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 80:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_x_8 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 69:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_x_8 <= io_matrixIn_8_re; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 80:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_x_9 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 69:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_x_9 <= io_matrixIn_9_re; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 80:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_y_0 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 70:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_y_0 <= io_matrixIn_0_im; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 81:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_y_1 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 70:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_y_1 <= io_matrixIn_1_im; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 81:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_y_2 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 70:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_y_2 <= io_matrixIn_2_im; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 81:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_y_3 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 70:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_y_3 <= io_matrixIn_3_im; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 81:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_y_4 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 70:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_y_4 <= io_matrixIn_4_im; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 81:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_y_5 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 70:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_y_5 <= io_matrixIn_5_im; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 81:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_y_6 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 70:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_y_6 <= io_matrixIn_6_im; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 81:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_y_7 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 70:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_y_7 <= io_matrixIn_7_im; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 81:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_y_8 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 70:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_y_8 <= io_matrixIn_8_im; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 81:16]
    end
    if (io_reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 67:18]
      reg_y_9 <= 64'sh0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 70:16]
    end else if (io_ready) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 77:24]
      reg_y_9 <= io_matrixIn_9_im; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 81:16]
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_0 <= _GEN_23;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      if (lower_tri_mat_inv_unit_io_valid) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 94:43]
        reg_x_inv_0 <= lower_tri_mat_inv_unit_io_matrixOut_0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 97:17]
      end else begin
        reg_x_inv_0 <= _GEN_23;
      end
    end else begin
      reg_x_inv_0 <= _GEN_23;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_1 <= _GEN_29;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      if (lower_tri_mat_inv_unit_io_valid) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 94:43]
        reg_x_inv_1 <= lower_tri_mat_inv_unit_io_matrixOut_1; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 97:17]
      end else begin
        reg_x_inv_1 <= _GEN_29;
      end
    end else begin
      reg_x_inv_1 <= _GEN_29;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_2 <= _GEN_35;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      if (lower_tri_mat_inv_unit_io_valid) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 94:43]
        reg_x_inv_2 <= lower_tri_mat_inv_unit_io_matrixOut_2; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 97:17]
      end else begin
        reg_x_inv_2 <= _GEN_35;
      end
    end else begin
      reg_x_inv_2 <= _GEN_35;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_3 <= _GEN_41;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      if (lower_tri_mat_inv_unit_io_valid) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 94:43]
        reg_x_inv_3 <= lower_tri_mat_inv_unit_io_matrixOut_3; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 97:17]
      end else begin
        reg_x_inv_3 <= _GEN_41;
      end
    end else begin
      reg_x_inv_3 <= _GEN_41;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_4 <= _GEN_47;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      if (lower_tri_mat_inv_unit_io_valid) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 94:43]
        reg_x_inv_4 <= lower_tri_mat_inv_unit_io_matrixOut_4; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 97:17]
      end else begin
        reg_x_inv_4 <= _GEN_47;
      end
    end else begin
      reg_x_inv_4 <= _GEN_47;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_5 <= _GEN_53;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      if (lower_tri_mat_inv_unit_io_valid) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 94:43]
        reg_x_inv_5 <= lower_tri_mat_inv_unit_io_matrixOut_5; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 97:17]
      end else begin
        reg_x_inv_5 <= _GEN_53;
      end
    end else begin
      reg_x_inv_5 <= _GEN_53;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_6 <= _GEN_59;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      if (lower_tri_mat_inv_unit_io_valid) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 94:43]
        reg_x_inv_6 <= lower_tri_mat_inv_unit_io_matrixOut_6; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 97:17]
      end else begin
        reg_x_inv_6 <= _GEN_59;
      end
    end else begin
      reg_x_inv_6 <= _GEN_59;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_7 <= _GEN_65;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      if (lower_tri_mat_inv_unit_io_valid) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 94:43]
        reg_x_inv_7 <= lower_tri_mat_inv_unit_io_matrixOut_7; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 97:17]
      end else begin
        reg_x_inv_7 <= _GEN_65;
      end
    end else begin
      reg_x_inv_7 <= _GEN_65;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_8 <= _GEN_71;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      if (lower_tri_mat_inv_unit_io_valid) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 94:43]
        reg_x_inv_8 <= lower_tri_mat_inv_unit_io_matrixOut_8; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 97:17]
      end else begin
        reg_x_inv_8 <= _GEN_71;
      end
    end else begin
      reg_x_inv_8 <= _GEN_71;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_9 <= _GEN_77;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      if (lower_tri_mat_inv_unit_io_valid) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 94:43]
        reg_x_inv_9 <= lower_tri_mat_inv_unit_io_matrixOut_9; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 97:17]
      end else begin
        reg_x_inv_9 <= _GEN_77;
      end
    end else begin
      reg_x_inv_9 <= _GEN_77;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_y_0 <= _GEN_24;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_x_inv_y_0 <= _GEN_24;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_x_inv_y_0 <= _GEN_24;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_x_inv_y_0 <= _GEN_94;
    end else begin
      reg_x_inv_y_0 <= _GEN_24;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_y_1 <= _GEN_30;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_x_inv_y_1 <= _GEN_30;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_x_inv_y_1 <= _GEN_30;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_x_inv_y_1 <= _GEN_95;
    end else begin
      reg_x_inv_y_1 <= _GEN_30;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_y_2 <= _GEN_36;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_x_inv_y_2 <= _GEN_36;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_x_inv_y_2 <= _GEN_36;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_x_inv_y_2 <= _GEN_96;
    end else begin
      reg_x_inv_y_2 <= _GEN_36;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_y_3 <= _GEN_42;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_x_inv_y_3 <= _GEN_42;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_x_inv_y_3 <= _GEN_42;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_x_inv_y_3 <= _GEN_97;
    end else begin
      reg_x_inv_y_3 <= _GEN_42;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_y_4 <= _GEN_48;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_x_inv_y_4 <= _GEN_48;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_x_inv_y_4 <= _GEN_48;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_x_inv_y_4 <= _GEN_98;
    end else begin
      reg_x_inv_y_4 <= _GEN_48;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_y_5 <= _GEN_54;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_x_inv_y_5 <= _GEN_54;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_x_inv_y_5 <= _GEN_54;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_x_inv_y_5 <= _GEN_99;
    end else begin
      reg_x_inv_y_5 <= _GEN_54;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_y_6 <= _GEN_60;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_x_inv_y_6 <= _GEN_60;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_x_inv_y_6 <= _GEN_60;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_x_inv_y_6 <= _GEN_100;
    end else begin
      reg_x_inv_y_6 <= _GEN_60;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_y_7 <= _GEN_66;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_x_inv_y_7 <= _GEN_66;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_x_inv_y_7 <= _GEN_66;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_x_inv_y_7 <= _GEN_101;
    end else begin
      reg_x_inv_y_7 <= _GEN_66;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_y_8 <= _GEN_72;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_x_inv_y_8 <= _GEN_72;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_x_inv_y_8 <= _GEN_72;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_x_inv_y_8 <= _GEN_102;
    end else begin
      reg_x_inv_y_8 <= _GEN_72;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_x_inv_y_9 <= _GEN_78;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_x_inv_y_9 <= _GEN_78;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_x_inv_y_9 <= _GEN_78;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_x_inv_y_9 <= _GEN_103;
    end else begin
      reg_x_inv_y_9 <= _GEN_78;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_u_0 <= _GEN_25;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_u_0 <= _GEN_25;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_u_0 <= _GEN_25;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_u_0 <= _GEN_25;
    end else begin
      reg_u_0 <= _GEN_357;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_u_1 <= _GEN_31;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_u_1 <= _GEN_31;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_u_1 <= _GEN_31;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_u_1 <= _GEN_31;
    end else begin
      reg_u_1 <= _GEN_358;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_u_2 <= _GEN_37;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_u_2 <= _GEN_37;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_u_2 <= _GEN_37;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_u_2 <= _GEN_37;
    end else begin
      reg_u_2 <= _GEN_359;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_u_3 <= _GEN_43;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_u_3 <= _GEN_43;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_u_3 <= _GEN_43;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_u_3 <= _GEN_43;
    end else begin
      reg_u_3 <= _GEN_360;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_u_4 <= _GEN_49;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_u_4 <= _GEN_49;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_u_4 <= _GEN_49;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_u_4 <= _GEN_49;
    end else begin
      reg_u_4 <= _GEN_361;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_u_5 <= _GEN_55;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_u_5 <= _GEN_55;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_u_5 <= _GEN_55;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_u_5 <= _GEN_55;
    end else begin
      reg_u_5 <= _GEN_362;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_u_6 <= _GEN_61;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_u_6 <= _GEN_61;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_u_6 <= _GEN_61;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_u_6 <= _GEN_61;
    end else begin
      reg_u_6 <= _GEN_363;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_u_7 <= _GEN_67;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_u_7 <= _GEN_67;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_u_7 <= _GEN_67;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_u_7 <= _GEN_67;
    end else begin
      reg_u_7 <= _GEN_364;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_u_8 <= _GEN_73;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_u_8 <= _GEN_73;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_u_8 <= _GEN_73;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_u_8 <= _GEN_73;
    end else begin
      reg_u_8 <= _GEN_365;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_u_9 <= _GEN_79;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_u_9 <= _GEN_79;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_u_9 <= _GEN_79;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_u_9 <= _GEN_79;
    end else begin
      reg_u_9 <= _GEN_366;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_v_0 <= _GEN_26;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_v_0 <= _GEN_26;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_v_0 <= _GEN_26;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_v_0 <= _GEN_26;
    end else begin
      reg_v_0 <= _GEN_378;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_v_1 <= _GEN_32;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_v_1 <= _GEN_32;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_v_1 <= _GEN_32;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_v_1 <= _GEN_32;
    end else begin
      reg_v_1 <= _GEN_379;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_v_2 <= _GEN_38;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_v_2 <= _GEN_38;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_v_2 <= _GEN_38;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_v_2 <= _GEN_38;
    end else begin
      reg_v_2 <= _GEN_380;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_v_3 <= _GEN_44;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_v_3 <= _GEN_44;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_v_3 <= _GEN_44;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_v_3 <= _GEN_44;
    end else begin
      reg_v_3 <= _GEN_381;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_v_4 <= _GEN_50;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_v_4 <= _GEN_50;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_v_4 <= _GEN_50;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_v_4 <= _GEN_50;
    end else begin
      reg_v_4 <= _GEN_382;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_v_5 <= _GEN_56;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_v_5 <= _GEN_56;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_v_5 <= _GEN_56;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_v_5 <= _GEN_56;
    end else begin
      reg_v_5 <= _GEN_383;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_v_6 <= _GEN_62;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_v_6 <= _GEN_62;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_v_6 <= _GEN_62;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_v_6 <= _GEN_62;
    end else begin
      reg_v_6 <= _GEN_384;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_v_7 <= _GEN_68;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_v_7 <= _GEN_68;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_v_7 <= _GEN_68;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_v_7 <= _GEN_68;
    end else begin
      reg_v_7 <= _GEN_385;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_v_8 <= _GEN_74;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_v_8 <= _GEN_74;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_v_8 <= _GEN_74;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_v_8 <= _GEN_74;
    end else begin
      reg_v_8 <= _GEN_386;
    end
    if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_v_9 <= _GEN_80;
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      reg_v_9 <= _GEN_80;
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_v_9 <= _GEN_80;
    end else if (reg_step_status == 4'h4) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 113:39]
      reg_v_9 <= _GEN_80;
    end else begin
      reg_v_9 <= _GEN_387;
    end
    if (reset) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 42:38]
      reg_step_status <= 4'h0; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 42:38]
    end else if (reg_step_status == 4'h1) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 86:33]
      reg_step_status <= _reg_step_status_T_1; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 90:21]
    end else if (reg_step_status == 4'h2) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 91:39]
      if (lower_tri_mat_inv_unit_io_valid) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 94:43]
        reg_step_status <= _reg_step_status_T_1; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 96:23]
      end else begin
        reg_step_status <= _GEN_81;
      end
    end else if (reg_step_status == 4'h3) begin // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 99:39]
      reg_step_status <= _reg_step_status_T_1; // @[Lower_Triangular_Matrix_Inversion_Complex_V1.scala 112:21]
    end else begin
      reg_step_status <= _GEN_389;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  reg_x_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  reg_x_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  reg_x_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  reg_x_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  reg_x_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  reg_x_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  reg_x_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  reg_x_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  reg_x_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  reg_x_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  reg_y_0 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  reg_y_1 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  reg_y_2 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  reg_y_3 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  reg_y_4 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  reg_y_5 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  reg_y_6 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  reg_y_7 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  reg_y_8 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  reg_y_9 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  reg_x_inv_0 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  reg_x_inv_1 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  reg_x_inv_2 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  reg_x_inv_3 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  reg_x_inv_4 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  reg_x_inv_5 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  reg_x_inv_6 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  reg_x_inv_7 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  reg_x_inv_8 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  reg_x_inv_9 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  reg_x_inv_y_0 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  reg_x_inv_y_1 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  reg_x_inv_y_2 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  reg_x_inv_y_3 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  reg_x_inv_y_4 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  reg_x_inv_y_5 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  reg_x_inv_y_6 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  reg_x_inv_y_7 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  reg_x_inv_y_8 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  reg_x_inv_y_9 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  reg_u_0 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  reg_u_1 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  reg_u_2 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  reg_u_3 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  reg_u_4 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  reg_u_5 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  reg_u_6 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  reg_u_7 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  reg_u_8 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  reg_u_9 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  reg_v_0 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  reg_v_1 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  reg_v_2 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  reg_v_3 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  reg_v_4 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  reg_v_5 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  reg_v_6 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  reg_v_7 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  reg_v_8 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  reg_v_9 = _RAND_59[63:0];
  _RAND_60 = {1{`RANDOM}};
  reg_step_status = _RAND_60[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module matrix_mul_v1_2(
  input         clock,
  input         io_reset,
  input         io_ready,
  input  [63:0] io_matrixA_0_re,
  input  [63:0] io_matrixA_0_im,
  input  [63:0] io_matrixA_1_re,
  input  [63:0] io_matrixA_1_im,
  input  [63:0] io_matrixA_2_re,
  input  [63:0] io_matrixA_2_im,
  input  [63:0] io_matrixA_3_re,
  input  [63:0] io_matrixA_3_im,
  input  [63:0] io_matrixA_5_re,
  input  [63:0] io_matrixA_5_im,
  input  [63:0] io_matrixA_6_re,
  input  [63:0] io_matrixA_6_im,
  input  [63:0] io_matrixA_7_re,
  input  [63:0] io_matrixA_7_im,
  input  [63:0] io_matrixA_10_re,
  input  [63:0] io_matrixA_10_im,
  input  [63:0] io_matrixA_11_re,
  input  [63:0] io_matrixA_11_im,
  input  [63:0] io_matrixA_15_re,
  input  [63:0] io_matrixA_15_im,
  input  [63:0] io_matrixB_0_re,
  input  [63:0] io_matrixB_0_im,
  input  [63:0] io_matrixB_4_re,
  input  [63:0] io_matrixB_4_im,
  input  [63:0] io_matrixB_5_re,
  input  [63:0] io_matrixB_5_im,
  input  [63:0] io_matrixB_8_re,
  input  [63:0] io_matrixB_8_im,
  input  [63:0] io_matrixB_9_re,
  input  [63:0] io_matrixB_9_im,
  input  [63:0] io_matrixB_10_re,
  input  [63:0] io_matrixB_10_im,
  input  [63:0] io_matrixB_12_re,
  input  [63:0] io_matrixB_12_im,
  input  [63:0] io_matrixB_13_re,
  input  [63:0] io_matrixB_13_im,
  input  [63:0] io_matrixB_14_re,
  input  [63:0] io_matrixB_14_im,
  input  [63:0] io_matrixB_15_re,
  input  [63:0] io_matrixB_15_im,
  output [63:0] io_matrixC_0_re,
  output [63:0] io_matrixC_0_im,
  output [63:0] io_matrixC_1_re,
  output [63:0] io_matrixC_1_im,
  output [63:0] io_matrixC_2_re,
  output [63:0] io_matrixC_2_im,
  output [63:0] io_matrixC_3_re,
  output [63:0] io_matrixC_3_im,
  output [63:0] io_matrixC_4_re,
  output [63:0] io_matrixC_4_im,
  output [63:0] io_matrixC_5_re,
  output [63:0] io_matrixC_5_im,
  output [63:0] io_matrixC_6_re,
  output [63:0] io_matrixC_6_im,
  output [63:0] io_matrixC_7_re,
  output [63:0] io_matrixC_7_im,
  output [63:0] io_matrixC_8_re,
  output [63:0] io_matrixC_8_im,
  output [63:0] io_matrixC_9_re,
  output [63:0] io_matrixC_9_im,
  output [63:0] io_matrixC_10_re,
  output [63:0] io_matrixC_10_im,
  output [63:0] io_matrixC_11_re,
  output [63:0] io_matrixC_11_im,
  output [63:0] io_matrixC_12_re,
  output [63:0] io_matrixC_12_im,
  output [63:0] io_matrixC_13_re,
  output [63:0] io_matrixC_13_im,
  output [63:0] io_matrixC_14_re,
  output [63:0] io_matrixC_14_im,
  output [63:0] io_matrixC_15_re,
  output [63:0] io_matrixC_15_im,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [31:0] _RAND_40;
`endif // RANDOMIZE_REG_INIT
  wire  PE_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_1_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_1_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_2_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_2_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_3_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_3_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_4_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_4_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_4_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_5_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_5_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_5_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_6_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_6_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_6_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_7_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_7_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_7_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_8_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_8_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_8_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_9_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_9_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_9_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_10_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_10_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_10_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_11_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_11_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_11_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_12_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_12_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_12_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_13_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_13_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_13_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_14_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_14_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_14_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_15_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_15_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_15_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  reg [63:0] regsA_0_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_0_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_1_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_1_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_2_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_2_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_3_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_3_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_5_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_5_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_6_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_6_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_7_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_7_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_10_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_10_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_11_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_11_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_15_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_15_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsB_0_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_0_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_4_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_4_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_5_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_5_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_8_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_8_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_9_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_9_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_10_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_10_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_12_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_12_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_13_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_13_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_14_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_14_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_15_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_15_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [4:0] input_point; // @[Matrix_Mul_V1.scala 84:30]
  wire [4:0] _input_point_T_1 = input_point + 5'h1; // @[Matrix_Mul_V1.scala 116:32]
  wire  _T = input_point < 5'h7; // @[Matrix_Mul_V1.scala 145:20]
  wire [3:0] _T_1 = 1'h0 * 3'h7; // @[Matrix_Mul_V1.scala 148:44]
  wire [4:0] _GEN_597 = {{1'd0}, _T_1}; // @[Matrix_Mul_V1.scala 148:60]
  wire [4:0] _T_3 = _GEN_597 + input_point; // @[Matrix_Mul_V1.scala 148:60]
  wire [63:0] _GEN_133 = 5'h1 == _T_3 ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_134 = 5'h2 == _T_3 ? $signed(regsA_2_im) : $signed(_GEN_133); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_135 = 5'h3 == _T_3 ? $signed(regsA_3_im) : $signed(_GEN_134); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_136 = 5'h4 == _T_3 ? $signed(64'sh0) : $signed(_GEN_135); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_137 = 5'h5 == _T_3 ? $signed(64'sh0) : $signed(_GEN_136); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_138 = 5'h6 == _T_3 ? $signed(64'sh0) : $signed(_GEN_137); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_139 = 5'h7 == _T_3 ? $signed(64'sh0) : $signed(_GEN_138); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_140 = 5'h8 == _T_3 ? $signed(64'sh0) : $signed(_GEN_139); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_141 = 5'h9 == _T_3 ? $signed(regsA_5_im) : $signed(_GEN_140); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_142 = 5'ha == _T_3 ? $signed(regsA_6_im) : $signed(_GEN_141); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_143 = 5'hb == _T_3 ? $signed(regsA_7_im) : $signed(_GEN_142); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_144 = 5'hc == _T_3 ? $signed(64'sh0) : $signed(_GEN_143); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_145 = 5'hd == _T_3 ? $signed(64'sh0) : $signed(_GEN_144); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_146 = 5'he == _T_3 ? $signed(64'sh0) : $signed(_GEN_145); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_147 = 5'hf == _T_3 ? $signed(64'sh0) : $signed(_GEN_146); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_148 = 5'h10 == _T_3 ? $signed(64'sh0) : $signed(_GEN_147); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_149 = 5'h11 == _T_3 ? $signed(64'sh0) : $signed(_GEN_148); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_150 = 5'h12 == _T_3 ? $signed(regsA_10_im) : $signed(_GEN_149); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_151 = 5'h13 == _T_3 ? $signed(regsA_11_im) : $signed(_GEN_150); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_152 = 5'h14 == _T_3 ? $signed(64'sh0) : $signed(_GEN_151); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_153 = 5'h15 == _T_3 ? $signed(64'sh0) : $signed(_GEN_152); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_154 = 5'h16 == _T_3 ? $signed(64'sh0) : $signed(_GEN_153); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_155 = 5'h17 == _T_3 ? $signed(64'sh0) : $signed(_GEN_154); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_156 = 5'h18 == _T_3 ? $signed(64'sh0) : $signed(_GEN_155); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_157 = 5'h19 == _T_3 ? $signed(64'sh0) : $signed(_GEN_156); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_158 = 5'h1a == _T_3 ? $signed(64'sh0) : $signed(_GEN_157); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_159 = 5'h1b == _T_3 ? $signed(regsA_15_im) : $signed(_GEN_158); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_161 = 5'h1 == _T_3 ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_162 = 5'h2 == _T_3 ? $signed(regsA_2_re) : $signed(_GEN_161); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_163 = 5'h3 == _T_3 ? $signed(regsA_3_re) : $signed(_GEN_162); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_164 = 5'h4 == _T_3 ? $signed(64'sh0) : $signed(_GEN_163); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_165 = 5'h5 == _T_3 ? $signed(64'sh0) : $signed(_GEN_164); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_166 = 5'h6 == _T_3 ? $signed(64'sh0) : $signed(_GEN_165); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_167 = 5'h7 == _T_3 ? $signed(64'sh0) : $signed(_GEN_166); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_168 = 5'h8 == _T_3 ? $signed(64'sh0) : $signed(_GEN_167); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_169 = 5'h9 == _T_3 ? $signed(regsA_5_re) : $signed(_GEN_168); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_170 = 5'ha == _T_3 ? $signed(regsA_6_re) : $signed(_GEN_169); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_171 = 5'hb == _T_3 ? $signed(regsA_7_re) : $signed(_GEN_170); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_172 = 5'hc == _T_3 ? $signed(64'sh0) : $signed(_GEN_171); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_173 = 5'hd == _T_3 ? $signed(64'sh0) : $signed(_GEN_172); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_174 = 5'he == _T_3 ? $signed(64'sh0) : $signed(_GEN_173); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_175 = 5'hf == _T_3 ? $signed(64'sh0) : $signed(_GEN_174); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_176 = 5'h10 == _T_3 ? $signed(64'sh0) : $signed(_GEN_175); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_177 = 5'h11 == _T_3 ? $signed(64'sh0) : $signed(_GEN_176); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_178 = 5'h12 == _T_3 ? $signed(regsA_10_re) : $signed(_GEN_177); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_179 = 5'h13 == _T_3 ? $signed(regsA_11_re) : $signed(_GEN_178); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_180 = 5'h14 == _T_3 ? $signed(64'sh0) : $signed(_GEN_179); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_181 = 5'h15 == _T_3 ? $signed(64'sh0) : $signed(_GEN_180); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_182 = 5'h16 == _T_3 ? $signed(64'sh0) : $signed(_GEN_181); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_183 = 5'h17 == _T_3 ? $signed(64'sh0) : $signed(_GEN_182); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_184 = 5'h18 == _T_3 ? $signed(64'sh0) : $signed(_GEN_183); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_185 = 5'h19 == _T_3 ? $signed(64'sh0) : $signed(_GEN_184); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_186 = 5'h1a == _T_3 ? $signed(64'sh0) : $signed(_GEN_185); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_187 = 5'h1b == _T_3 ? $signed(regsA_15_re) : $signed(_GEN_186); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [3:0] _T_4 = 1'h1 * 3'h7; // @[Matrix_Mul_V1.scala 148:44]
  wire [4:0] _GEN_598 = {{1'd0}, _T_4}; // @[Matrix_Mul_V1.scala 148:60]
  wire [4:0] _T_6 = _GEN_598 + input_point; // @[Matrix_Mul_V1.scala 148:60]
  wire [63:0] _GEN_189 = 5'h1 == _T_6 ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_190 = 5'h2 == _T_6 ? $signed(regsA_2_im) : $signed(_GEN_189); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_191 = 5'h3 == _T_6 ? $signed(regsA_3_im) : $signed(_GEN_190); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_192 = 5'h4 == _T_6 ? $signed(64'sh0) : $signed(_GEN_191); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_193 = 5'h5 == _T_6 ? $signed(64'sh0) : $signed(_GEN_192); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_194 = 5'h6 == _T_6 ? $signed(64'sh0) : $signed(_GEN_193); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_195 = 5'h7 == _T_6 ? $signed(64'sh0) : $signed(_GEN_194); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_196 = 5'h8 == _T_6 ? $signed(64'sh0) : $signed(_GEN_195); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_197 = 5'h9 == _T_6 ? $signed(regsA_5_im) : $signed(_GEN_196); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_198 = 5'ha == _T_6 ? $signed(regsA_6_im) : $signed(_GEN_197); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_199 = 5'hb == _T_6 ? $signed(regsA_7_im) : $signed(_GEN_198); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_200 = 5'hc == _T_6 ? $signed(64'sh0) : $signed(_GEN_199); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_201 = 5'hd == _T_6 ? $signed(64'sh0) : $signed(_GEN_200); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_202 = 5'he == _T_6 ? $signed(64'sh0) : $signed(_GEN_201); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_203 = 5'hf == _T_6 ? $signed(64'sh0) : $signed(_GEN_202); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_204 = 5'h10 == _T_6 ? $signed(64'sh0) : $signed(_GEN_203); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_205 = 5'h11 == _T_6 ? $signed(64'sh0) : $signed(_GEN_204); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_206 = 5'h12 == _T_6 ? $signed(regsA_10_im) : $signed(_GEN_205); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_207 = 5'h13 == _T_6 ? $signed(regsA_11_im) : $signed(_GEN_206); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_208 = 5'h14 == _T_6 ? $signed(64'sh0) : $signed(_GEN_207); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_209 = 5'h15 == _T_6 ? $signed(64'sh0) : $signed(_GEN_208); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_210 = 5'h16 == _T_6 ? $signed(64'sh0) : $signed(_GEN_209); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_211 = 5'h17 == _T_6 ? $signed(64'sh0) : $signed(_GEN_210); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_212 = 5'h18 == _T_6 ? $signed(64'sh0) : $signed(_GEN_211); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_213 = 5'h19 == _T_6 ? $signed(64'sh0) : $signed(_GEN_212); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_214 = 5'h1a == _T_6 ? $signed(64'sh0) : $signed(_GEN_213); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_215 = 5'h1b == _T_6 ? $signed(regsA_15_im) : $signed(_GEN_214); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_217 = 5'h1 == _T_6 ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_218 = 5'h2 == _T_6 ? $signed(regsA_2_re) : $signed(_GEN_217); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_219 = 5'h3 == _T_6 ? $signed(regsA_3_re) : $signed(_GEN_218); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_220 = 5'h4 == _T_6 ? $signed(64'sh0) : $signed(_GEN_219); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_221 = 5'h5 == _T_6 ? $signed(64'sh0) : $signed(_GEN_220); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_222 = 5'h6 == _T_6 ? $signed(64'sh0) : $signed(_GEN_221); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_223 = 5'h7 == _T_6 ? $signed(64'sh0) : $signed(_GEN_222); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_224 = 5'h8 == _T_6 ? $signed(64'sh0) : $signed(_GEN_223); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_225 = 5'h9 == _T_6 ? $signed(regsA_5_re) : $signed(_GEN_224); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_226 = 5'ha == _T_6 ? $signed(regsA_6_re) : $signed(_GEN_225); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_227 = 5'hb == _T_6 ? $signed(regsA_7_re) : $signed(_GEN_226); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_228 = 5'hc == _T_6 ? $signed(64'sh0) : $signed(_GEN_227); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_229 = 5'hd == _T_6 ? $signed(64'sh0) : $signed(_GEN_228); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_230 = 5'he == _T_6 ? $signed(64'sh0) : $signed(_GEN_229); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_231 = 5'hf == _T_6 ? $signed(64'sh0) : $signed(_GEN_230); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_232 = 5'h10 == _T_6 ? $signed(64'sh0) : $signed(_GEN_231); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_233 = 5'h11 == _T_6 ? $signed(64'sh0) : $signed(_GEN_232); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_234 = 5'h12 == _T_6 ? $signed(regsA_10_re) : $signed(_GEN_233); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_235 = 5'h13 == _T_6 ? $signed(regsA_11_re) : $signed(_GEN_234); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_236 = 5'h14 == _T_6 ? $signed(64'sh0) : $signed(_GEN_235); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_237 = 5'h15 == _T_6 ? $signed(64'sh0) : $signed(_GEN_236); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_238 = 5'h16 == _T_6 ? $signed(64'sh0) : $signed(_GEN_237); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_239 = 5'h17 == _T_6 ? $signed(64'sh0) : $signed(_GEN_238); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_240 = 5'h18 == _T_6 ? $signed(64'sh0) : $signed(_GEN_239); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_241 = 5'h19 == _T_6 ? $signed(64'sh0) : $signed(_GEN_240); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_242 = 5'h1a == _T_6 ? $signed(64'sh0) : $signed(_GEN_241); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_243 = 5'h1b == _T_6 ? $signed(regsA_15_re) : $signed(_GEN_242); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [4:0] _T_7 = 2'h2 * 3'h7; // @[Matrix_Mul_V1.scala 148:44]
  wire [4:0] _T_9 = _T_7 + input_point; // @[Matrix_Mul_V1.scala 148:60]
  wire [63:0] _GEN_245 = 5'h1 == _T_9 ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_246 = 5'h2 == _T_9 ? $signed(regsA_2_im) : $signed(_GEN_245); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_247 = 5'h3 == _T_9 ? $signed(regsA_3_im) : $signed(_GEN_246); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_248 = 5'h4 == _T_9 ? $signed(64'sh0) : $signed(_GEN_247); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_249 = 5'h5 == _T_9 ? $signed(64'sh0) : $signed(_GEN_248); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_250 = 5'h6 == _T_9 ? $signed(64'sh0) : $signed(_GEN_249); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_251 = 5'h7 == _T_9 ? $signed(64'sh0) : $signed(_GEN_250); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_252 = 5'h8 == _T_9 ? $signed(64'sh0) : $signed(_GEN_251); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_253 = 5'h9 == _T_9 ? $signed(regsA_5_im) : $signed(_GEN_252); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_254 = 5'ha == _T_9 ? $signed(regsA_6_im) : $signed(_GEN_253); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_255 = 5'hb == _T_9 ? $signed(regsA_7_im) : $signed(_GEN_254); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_256 = 5'hc == _T_9 ? $signed(64'sh0) : $signed(_GEN_255); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_257 = 5'hd == _T_9 ? $signed(64'sh0) : $signed(_GEN_256); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_258 = 5'he == _T_9 ? $signed(64'sh0) : $signed(_GEN_257); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_259 = 5'hf == _T_9 ? $signed(64'sh0) : $signed(_GEN_258); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_260 = 5'h10 == _T_9 ? $signed(64'sh0) : $signed(_GEN_259); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_261 = 5'h11 == _T_9 ? $signed(64'sh0) : $signed(_GEN_260); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_262 = 5'h12 == _T_9 ? $signed(regsA_10_im) : $signed(_GEN_261); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_263 = 5'h13 == _T_9 ? $signed(regsA_11_im) : $signed(_GEN_262); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_264 = 5'h14 == _T_9 ? $signed(64'sh0) : $signed(_GEN_263); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_265 = 5'h15 == _T_9 ? $signed(64'sh0) : $signed(_GEN_264); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_266 = 5'h16 == _T_9 ? $signed(64'sh0) : $signed(_GEN_265); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_267 = 5'h17 == _T_9 ? $signed(64'sh0) : $signed(_GEN_266); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_268 = 5'h18 == _T_9 ? $signed(64'sh0) : $signed(_GEN_267); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_269 = 5'h19 == _T_9 ? $signed(64'sh0) : $signed(_GEN_268); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_270 = 5'h1a == _T_9 ? $signed(64'sh0) : $signed(_GEN_269); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_271 = 5'h1b == _T_9 ? $signed(regsA_15_im) : $signed(_GEN_270); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_273 = 5'h1 == _T_9 ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_274 = 5'h2 == _T_9 ? $signed(regsA_2_re) : $signed(_GEN_273); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_275 = 5'h3 == _T_9 ? $signed(regsA_3_re) : $signed(_GEN_274); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_276 = 5'h4 == _T_9 ? $signed(64'sh0) : $signed(_GEN_275); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_277 = 5'h5 == _T_9 ? $signed(64'sh0) : $signed(_GEN_276); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_278 = 5'h6 == _T_9 ? $signed(64'sh0) : $signed(_GEN_277); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_279 = 5'h7 == _T_9 ? $signed(64'sh0) : $signed(_GEN_278); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_280 = 5'h8 == _T_9 ? $signed(64'sh0) : $signed(_GEN_279); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_281 = 5'h9 == _T_9 ? $signed(regsA_5_re) : $signed(_GEN_280); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_282 = 5'ha == _T_9 ? $signed(regsA_6_re) : $signed(_GEN_281); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_283 = 5'hb == _T_9 ? $signed(regsA_7_re) : $signed(_GEN_282); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_284 = 5'hc == _T_9 ? $signed(64'sh0) : $signed(_GEN_283); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_285 = 5'hd == _T_9 ? $signed(64'sh0) : $signed(_GEN_284); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_286 = 5'he == _T_9 ? $signed(64'sh0) : $signed(_GEN_285); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_287 = 5'hf == _T_9 ? $signed(64'sh0) : $signed(_GEN_286); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_288 = 5'h10 == _T_9 ? $signed(64'sh0) : $signed(_GEN_287); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_289 = 5'h11 == _T_9 ? $signed(64'sh0) : $signed(_GEN_288); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_290 = 5'h12 == _T_9 ? $signed(regsA_10_re) : $signed(_GEN_289); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_291 = 5'h13 == _T_9 ? $signed(regsA_11_re) : $signed(_GEN_290); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_292 = 5'h14 == _T_9 ? $signed(64'sh0) : $signed(_GEN_291); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_293 = 5'h15 == _T_9 ? $signed(64'sh0) : $signed(_GEN_292); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_294 = 5'h16 == _T_9 ? $signed(64'sh0) : $signed(_GEN_293); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_295 = 5'h17 == _T_9 ? $signed(64'sh0) : $signed(_GEN_294); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_296 = 5'h18 == _T_9 ? $signed(64'sh0) : $signed(_GEN_295); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_297 = 5'h19 == _T_9 ? $signed(64'sh0) : $signed(_GEN_296); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_298 = 5'h1a == _T_9 ? $signed(64'sh0) : $signed(_GEN_297); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_299 = 5'h1b == _T_9 ? $signed(regsA_15_re) : $signed(_GEN_298); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [4:0] _T_10 = 2'h3 * 3'h7; // @[Matrix_Mul_V1.scala 148:44]
  wire [4:0] _T_12 = _T_10 + input_point; // @[Matrix_Mul_V1.scala 148:60]
  wire [63:0] _GEN_301 = 5'h1 == _T_12 ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_302 = 5'h2 == _T_12 ? $signed(regsA_2_im) : $signed(_GEN_301); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_303 = 5'h3 == _T_12 ? $signed(regsA_3_im) : $signed(_GEN_302); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_304 = 5'h4 == _T_12 ? $signed(64'sh0) : $signed(_GEN_303); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_305 = 5'h5 == _T_12 ? $signed(64'sh0) : $signed(_GEN_304); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_306 = 5'h6 == _T_12 ? $signed(64'sh0) : $signed(_GEN_305); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_307 = 5'h7 == _T_12 ? $signed(64'sh0) : $signed(_GEN_306); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_308 = 5'h8 == _T_12 ? $signed(64'sh0) : $signed(_GEN_307); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_309 = 5'h9 == _T_12 ? $signed(regsA_5_im) : $signed(_GEN_308); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_310 = 5'ha == _T_12 ? $signed(regsA_6_im) : $signed(_GEN_309); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_311 = 5'hb == _T_12 ? $signed(regsA_7_im) : $signed(_GEN_310); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_312 = 5'hc == _T_12 ? $signed(64'sh0) : $signed(_GEN_311); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_313 = 5'hd == _T_12 ? $signed(64'sh0) : $signed(_GEN_312); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_314 = 5'he == _T_12 ? $signed(64'sh0) : $signed(_GEN_313); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_315 = 5'hf == _T_12 ? $signed(64'sh0) : $signed(_GEN_314); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_316 = 5'h10 == _T_12 ? $signed(64'sh0) : $signed(_GEN_315); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_317 = 5'h11 == _T_12 ? $signed(64'sh0) : $signed(_GEN_316); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_318 = 5'h12 == _T_12 ? $signed(regsA_10_im) : $signed(_GEN_317); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_319 = 5'h13 == _T_12 ? $signed(regsA_11_im) : $signed(_GEN_318); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_320 = 5'h14 == _T_12 ? $signed(64'sh0) : $signed(_GEN_319); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_321 = 5'h15 == _T_12 ? $signed(64'sh0) : $signed(_GEN_320); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_322 = 5'h16 == _T_12 ? $signed(64'sh0) : $signed(_GEN_321); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_323 = 5'h17 == _T_12 ? $signed(64'sh0) : $signed(_GEN_322); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_324 = 5'h18 == _T_12 ? $signed(64'sh0) : $signed(_GEN_323); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_325 = 5'h19 == _T_12 ? $signed(64'sh0) : $signed(_GEN_324); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_326 = 5'h1a == _T_12 ? $signed(64'sh0) : $signed(_GEN_325); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_327 = 5'h1b == _T_12 ? $signed(regsA_15_im) : $signed(_GEN_326); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_329 = 5'h1 == _T_12 ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_330 = 5'h2 == _T_12 ? $signed(regsA_2_re) : $signed(_GEN_329); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_331 = 5'h3 == _T_12 ? $signed(regsA_3_re) : $signed(_GEN_330); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_332 = 5'h4 == _T_12 ? $signed(64'sh0) : $signed(_GEN_331); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_333 = 5'h5 == _T_12 ? $signed(64'sh0) : $signed(_GEN_332); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_334 = 5'h6 == _T_12 ? $signed(64'sh0) : $signed(_GEN_333); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_335 = 5'h7 == _T_12 ? $signed(64'sh0) : $signed(_GEN_334); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_336 = 5'h8 == _T_12 ? $signed(64'sh0) : $signed(_GEN_335); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_337 = 5'h9 == _T_12 ? $signed(regsA_5_re) : $signed(_GEN_336); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_338 = 5'ha == _T_12 ? $signed(regsA_6_re) : $signed(_GEN_337); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_339 = 5'hb == _T_12 ? $signed(regsA_7_re) : $signed(_GEN_338); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_340 = 5'hc == _T_12 ? $signed(64'sh0) : $signed(_GEN_339); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_341 = 5'hd == _T_12 ? $signed(64'sh0) : $signed(_GEN_340); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_342 = 5'he == _T_12 ? $signed(64'sh0) : $signed(_GEN_341); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_343 = 5'hf == _T_12 ? $signed(64'sh0) : $signed(_GEN_342); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_344 = 5'h10 == _T_12 ? $signed(64'sh0) : $signed(_GEN_343); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_345 = 5'h11 == _T_12 ? $signed(64'sh0) : $signed(_GEN_344); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_346 = 5'h12 == _T_12 ? $signed(regsA_10_re) : $signed(_GEN_345); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_347 = 5'h13 == _T_12 ? $signed(regsA_11_re) : $signed(_GEN_346); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_348 = 5'h14 == _T_12 ? $signed(64'sh0) : $signed(_GEN_347); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_349 = 5'h15 == _T_12 ? $signed(64'sh0) : $signed(_GEN_348); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_350 = 5'h16 == _T_12 ? $signed(64'sh0) : $signed(_GEN_349); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_351 = 5'h17 == _T_12 ? $signed(64'sh0) : $signed(_GEN_350); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_352 = 5'h18 == _T_12 ? $signed(64'sh0) : $signed(_GEN_351); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_353 = 5'h19 == _T_12 ? $signed(64'sh0) : $signed(_GEN_352); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_354 = 5'h1a == _T_12 ? $signed(64'sh0) : $signed(_GEN_353); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_355 = 5'h1b == _T_12 ? $signed(regsA_15_re) : $signed(_GEN_354); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_365 = 5'h1 == _T_3 ? $signed(regsB_4_im) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_366 = 5'h2 == _T_3 ? $signed(regsB_8_im) : $signed(_GEN_365); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_367 = 5'h3 == _T_3 ? $signed(regsB_12_im) : $signed(_GEN_366); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_368 = 5'h4 == _T_3 ? $signed(64'sh0) : $signed(_GEN_367); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_369 = 5'h5 == _T_3 ? $signed(64'sh0) : $signed(_GEN_368); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_370 = 5'h6 == _T_3 ? $signed(64'sh0) : $signed(_GEN_369); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_371 = 5'h7 == _T_3 ? $signed(64'sh0) : $signed(_GEN_370); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_372 = 5'h8 == _T_3 ? $signed(64'sh0) : $signed(_GEN_371); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_373 = 5'h9 == _T_3 ? $signed(regsB_5_im) : $signed(_GEN_372); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_374 = 5'ha == _T_3 ? $signed(regsB_9_im) : $signed(_GEN_373); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_375 = 5'hb == _T_3 ? $signed(regsB_13_im) : $signed(_GEN_374); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_376 = 5'hc == _T_3 ? $signed(64'sh0) : $signed(_GEN_375); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_377 = 5'hd == _T_3 ? $signed(64'sh0) : $signed(_GEN_376); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_378 = 5'he == _T_3 ? $signed(64'sh0) : $signed(_GEN_377); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_379 = 5'hf == _T_3 ? $signed(64'sh0) : $signed(_GEN_378); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_380 = 5'h10 == _T_3 ? $signed(64'sh0) : $signed(_GEN_379); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_381 = 5'h11 == _T_3 ? $signed(64'sh0) : $signed(_GEN_380); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_382 = 5'h12 == _T_3 ? $signed(regsB_10_im) : $signed(_GEN_381); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_383 = 5'h13 == _T_3 ? $signed(regsB_14_im) : $signed(_GEN_382); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_384 = 5'h14 == _T_3 ? $signed(64'sh0) : $signed(_GEN_383); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_385 = 5'h15 == _T_3 ? $signed(64'sh0) : $signed(_GEN_384); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_386 = 5'h16 == _T_3 ? $signed(64'sh0) : $signed(_GEN_385); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_387 = 5'h17 == _T_3 ? $signed(64'sh0) : $signed(_GEN_386); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_388 = 5'h18 == _T_3 ? $signed(64'sh0) : $signed(_GEN_387); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_389 = 5'h19 == _T_3 ? $signed(64'sh0) : $signed(_GEN_388); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_390 = 5'h1a == _T_3 ? $signed(64'sh0) : $signed(_GEN_389); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_391 = 5'h1b == _T_3 ? $signed(regsB_15_im) : $signed(_GEN_390); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_393 = 5'h1 == _T_3 ? $signed(regsB_4_re) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_394 = 5'h2 == _T_3 ? $signed(regsB_8_re) : $signed(_GEN_393); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_395 = 5'h3 == _T_3 ? $signed(regsB_12_re) : $signed(_GEN_394); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_396 = 5'h4 == _T_3 ? $signed(64'sh0) : $signed(_GEN_395); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_397 = 5'h5 == _T_3 ? $signed(64'sh0) : $signed(_GEN_396); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_398 = 5'h6 == _T_3 ? $signed(64'sh0) : $signed(_GEN_397); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_399 = 5'h7 == _T_3 ? $signed(64'sh0) : $signed(_GEN_398); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_400 = 5'h8 == _T_3 ? $signed(64'sh0) : $signed(_GEN_399); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_401 = 5'h9 == _T_3 ? $signed(regsB_5_re) : $signed(_GEN_400); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_402 = 5'ha == _T_3 ? $signed(regsB_9_re) : $signed(_GEN_401); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_403 = 5'hb == _T_3 ? $signed(regsB_13_re) : $signed(_GEN_402); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_404 = 5'hc == _T_3 ? $signed(64'sh0) : $signed(_GEN_403); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_405 = 5'hd == _T_3 ? $signed(64'sh0) : $signed(_GEN_404); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_406 = 5'he == _T_3 ? $signed(64'sh0) : $signed(_GEN_405); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_407 = 5'hf == _T_3 ? $signed(64'sh0) : $signed(_GEN_406); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_408 = 5'h10 == _T_3 ? $signed(64'sh0) : $signed(_GEN_407); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_409 = 5'h11 == _T_3 ? $signed(64'sh0) : $signed(_GEN_408); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_410 = 5'h12 == _T_3 ? $signed(regsB_10_re) : $signed(_GEN_409); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_411 = 5'h13 == _T_3 ? $signed(regsB_14_re) : $signed(_GEN_410); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_412 = 5'h14 == _T_3 ? $signed(64'sh0) : $signed(_GEN_411); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_413 = 5'h15 == _T_3 ? $signed(64'sh0) : $signed(_GEN_412); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_414 = 5'h16 == _T_3 ? $signed(64'sh0) : $signed(_GEN_413); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_415 = 5'h17 == _T_3 ? $signed(64'sh0) : $signed(_GEN_414); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_416 = 5'h18 == _T_3 ? $signed(64'sh0) : $signed(_GEN_415); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_417 = 5'h19 == _T_3 ? $signed(64'sh0) : $signed(_GEN_416); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_418 = 5'h1a == _T_3 ? $signed(64'sh0) : $signed(_GEN_417); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_419 = 5'h1b == _T_3 ? $signed(regsB_15_re) : $signed(_GEN_418); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_421 = 5'h1 == _T_6 ? $signed(regsB_4_im) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_422 = 5'h2 == _T_6 ? $signed(regsB_8_im) : $signed(_GEN_421); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_423 = 5'h3 == _T_6 ? $signed(regsB_12_im) : $signed(_GEN_422); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_424 = 5'h4 == _T_6 ? $signed(64'sh0) : $signed(_GEN_423); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_425 = 5'h5 == _T_6 ? $signed(64'sh0) : $signed(_GEN_424); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_426 = 5'h6 == _T_6 ? $signed(64'sh0) : $signed(_GEN_425); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_427 = 5'h7 == _T_6 ? $signed(64'sh0) : $signed(_GEN_426); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_428 = 5'h8 == _T_6 ? $signed(64'sh0) : $signed(_GEN_427); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_429 = 5'h9 == _T_6 ? $signed(regsB_5_im) : $signed(_GEN_428); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_430 = 5'ha == _T_6 ? $signed(regsB_9_im) : $signed(_GEN_429); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_431 = 5'hb == _T_6 ? $signed(regsB_13_im) : $signed(_GEN_430); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_432 = 5'hc == _T_6 ? $signed(64'sh0) : $signed(_GEN_431); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_433 = 5'hd == _T_6 ? $signed(64'sh0) : $signed(_GEN_432); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_434 = 5'he == _T_6 ? $signed(64'sh0) : $signed(_GEN_433); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_435 = 5'hf == _T_6 ? $signed(64'sh0) : $signed(_GEN_434); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_436 = 5'h10 == _T_6 ? $signed(64'sh0) : $signed(_GEN_435); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_437 = 5'h11 == _T_6 ? $signed(64'sh0) : $signed(_GEN_436); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_438 = 5'h12 == _T_6 ? $signed(regsB_10_im) : $signed(_GEN_437); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_439 = 5'h13 == _T_6 ? $signed(regsB_14_im) : $signed(_GEN_438); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_440 = 5'h14 == _T_6 ? $signed(64'sh0) : $signed(_GEN_439); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_441 = 5'h15 == _T_6 ? $signed(64'sh0) : $signed(_GEN_440); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_442 = 5'h16 == _T_6 ? $signed(64'sh0) : $signed(_GEN_441); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_443 = 5'h17 == _T_6 ? $signed(64'sh0) : $signed(_GEN_442); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_444 = 5'h18 == _T_6 ? $signed(64'sh0) : $signed(_GEN_443); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_445 = 5'h19 == _T_6 ? $signed(64'sh0) : $signed(_GEN_444); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_446 = 5'h1a == _T_6 ? $signed(64'sh0) : $signed(_GEN_445); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_447 = 5'h1b == _T_6 ? $signed(regsB_15_im) : $signed(_GEN_446); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_449 = 5'h1 == _T_6 ? $signed(regsB_4_re) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_450 = 5'h2 == _T_6 ? $signed(regsB_8_re) : $signed(_GEN_449); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_451 = 5'h3 == _T_6 ? $signed(regsB_12_re) : $signed(_GEN_450); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_452 = 5'h4 == _T_6 ? $signed(64'sh0) : $signed(_GEN_451); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_453 = 5'h5 == _T_6 ? $signed(64'sh0) : $signed(_GEN_452); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_454 = 5'h6 == _T_6 ? $signed(64'sh0) : $signed(_GEN_453); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_455 = 5'h7 == _T_6 ? $signed(64'sh0) : $signed(_GEN_454); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_456 = 5'h8 == _T_6 ? $signed(64'sh0) : $signed(_GEN_455); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_457 = 5'h9 == _T_6 ? $signed(regsB_5_re) : $signed(_GEN_456); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_458 = 5'ha == _T_6 ? $signed(regsB_9_re) : $signed(_GEN_457); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_459 = 5'hb == _T_6 ? $signed(regsB_13_re) : $signed(_GEN_458); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_460 = 5'hc == _T_6 ? $signed(64'sh0) : $signed(_GEN_459); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_461 = 5'hd == _T_6 ? $signed(64'sh0) : $signed(_GEN_460); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_462 = 5'he == _T_6 ? $signed(64'sh0) : $signed(_GEN_461); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_463 = 5'hf == _T_6 ? $signed(64'sh0) : $signed(_GEN_462); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_464 = 5'h10 == _T_6 ? $signed(64'sh0) : $signed(_GEN_463); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_465 = 5'h11 == _T_6 ? $signed(64'sh0) : $signed(_GEN_464); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_466 = 5'h12 == _T_6 ? $signed(regsB_10_re) : $signed(_GEN_465); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_467 = 5'h13 == _T_6 ? $signed(regsB_14_re) : $signed(_GEN_466); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_468 = 5'h14 == _T_6 ? $signed(64'sh0) : $signed(_GEN_467); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_469 = 5'h15 == _T_6 ? $signed(64'sh0) : $signed(_GEN_468); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_470 = 5'h16 == _T_6 ? $signed(64'sh0) : $signed(_GEN_469); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_471 = 5'h17 == _T_6 ? $signed(64'sh0) : $signed(_GEN_470); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_472 = 5'h18 == _T_6 ? $signed(64'sh0) : $signed(_GEN_471); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_473 = 5'h19 == _T_6 ? $signed(64'sh0) : $signed(_GEN_472); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_474 = 5'h1a == _T_6 ? $signed(64'sh0) : $signed(_GEN_473); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_475 = 5'h1b == _T_6 ? $signed(regsB_15_re) : $signed(_GEN_474); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_477 = 5'h1 == _T_9 ? $signed(regsB_4_im) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_478 = 5'h2 == _T_9 ? $signed(regsB_8_im) : $signed(_GEN_477); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_479 = 5'h3 == _T_9 ? $signed(regsB_12_im) : $signed(_GEN_478); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_480 = 5'h4 == _T_9 ? $signed(64'sh0) : $signed(_GEN_479); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_481 = 5'h5 == _T_9 ? $signed(64'sh0) : $signed(_GEN_480); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_482 = 5'h6 == _T_9 ? $signed(64'sh0) : $signed(_GEN_481); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_483 = 5'h7 == _T_9 ? $signed(64'sh0) : $signed(_GEN_482); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_484 = 5'h8 == _T_9 ? $signed(64'sh0) : $signed(_GEN_483); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_485 = 5'h9 == _T_9 ? $signed(regsB_5_im) : $signed(_GEN_484); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_486 = 5'ha == _T_9 ? $signed(regsB_9_im) : $signed(_GEN_485); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_487 = 5'hb == _T_9 ? $signed(regsB_13_im) : $signed(_GEN_486); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_488 = 5'hc == _T_9 ? $signed(64'sh0) : $signed(_GEN_487); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_489 = 5'hd == _T_9 ? $signed(64'sh0) : $signed(_GEN_488); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_490 = 5'he == _T_9 ? $signed(64'sh0) : $signed(_GEN_489); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_491 = 5'hf == _T_9 ? $signed(64'sh0) : $signed(_GEN_490); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_492 = 5'h10 == _T_9 ? $signed(64'sh0) : $signed(_GEN_491); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_493 = 5'h11 == _T_9 ? $signed(64'sh0) : $signed(_GEN_492); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_494 = 5'h12 == _T_9 ? $signed(regsB_10_im) : $signed(_GEN_493); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_495 = 5'h13 == _T_9 ? $signed(regsB_14_im) : $signed(_GEN_494); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_496 = 5'h14 == _T_9 ? $signed(64'sh0) : $signed(_GEN_495); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_497 = 5'h15 == _T_9 ? $signed(64'sh0) : $signed(_GEN_496); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_498 = 5'h16 == _T_9 ? $signed(64'sh0) : $signed(_GEN_497); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_499 = 5'h17 == _T_9 ? $signed(64'sh0) : $signed(_GEN_498); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_500 = 5'h18 == _T_9 ? $signed(64'sh0) : $signed(_GEN_499); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_501 = 5'h19 == _T_9 ? $signed(64'sh0) : $signed(_GEN_500); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_502 = 5'h1a == _T_9 ? $signed(64'sh0) : $signed(_GEN_501); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_503 = 5'h1b == _T_9 ? $signed(regsB_15_im) : $signed(_GEN_502); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_505 = 5'h1 == _T_9 ? $signed(regsB_4_re) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_506 = 5'h2 == _T_9 ? $signed(regsB_8_re) : $signed(_GEN_505); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_507 = 5'h3 == _T_9 ? $signed(regsB_12_re) : $signed(_GEN_506); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_508 = 5'h4 == _T_9 ? $signed(64'sh0) : $signed(_GEN_507); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_509 = 5'h5 == _T_9 ? $signed(64'sh0) : $signed(_GEN_508); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_510 = 5'h6 == _T_9 ? $signed(64'sh0) : $signed(_GEN_509); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_511 = 5'h7 == _T_9 ? $signed(64'sh0) : $signed(_GEN_510); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_512 = 5'h8 == _T_9 ? $signed(64'sh0) : $signed(_GEN_511); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_513 = 5'h9 == _T_9 ? $signed(regsB_5_re) : $signed(_GEN_512); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_514 = 5'ha == _T_9 ? $signed(regsB_9_re) : $signed(_GEN_513); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_515 = 5'hb == _T_9 ? $signed(regsB_13_re) : $signed(_GEN_514); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_516 = 5'hc == _T_9 ? $signed(64'sh0) : $signed(_GEN_515); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_517 = 5'hd == _T_9 ? $signed(64'sh0) : $signed(_GEN_516); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_518 = 5'he == _T_9 ? $signed(64'sh0) : $signed(_GEN_517); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_519 = 5'hf == _T_9 ? $signed(64'sh0) : $signed(_GEN_518); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_520 = 5'h10 == _T_9 ? $signed(64'sh0) : $signed(_GEN_519); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_521 = 5'h11 == _T_9 ? $signed(64'sh0) : $signed(_GEN_520); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_522 = 5'h12 == _T_9 ? $signed(regsB_10_re) : $signed(_GEN_521); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_523 = 5'h13 == _T_9 ? $signed(regsB_14_re) : $signed(_GEN_522); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_524 = 5'h14 == _T_9 ? $signed(64'sh0) : $signed(_GEN_523); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_525 = 5'h15 == _T_9 ? $signed(64'sh0) : $signed(_GEN_524); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_526 = 5'h16 == _T_9 ? $signed(64'sh0) : $signed(_GEN_525); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_527 = 5'h17 == _T_9 ? $signed(64'sh0) : $signed(_GEN_526); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_528 = 5'h18 == _T_9 ? $signed(64'sh0) : $signed(_GEN_527); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_529 = 5'h19 == _T_9 ? $signed(64'sh0) : $signed(_GEN_528); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_530 = 5'h1a == _T_9 ? $signed(64'sh0) : $signed(_GEN_529); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_531 = 5'h1b == _T_9 ? $signed(regsB_15_re) : $signed(_GEN_530); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_533 = 5'h1 == _T_12 ? $signed(regsB_4_im) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_534 = 5'h2 == _T_12 ? $signed(regsB_8_im) : $signed(_GEN_533); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_535 = 5'h3 == _T_12 ? $signed(regsB_12_im) : $signed(_GEN_534); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_536 = 5'h4 == _T_12 ? $signed(64'sh0) : $signed(_GEN_535); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_537 = 5'h5 == _T_12 ? $signed(64'sh0) : $signed(_GEN_536); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_538 = 5'h6 == _T_12 ? $signed(64'sh0) : $signed(_GEN_537); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_539 = 5'h7 == _T_12 ? $signed(64'sh0) : $signed(_GEN_538); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_540 = 5'h8 == _T_12 ? $signed(64'sh0) : $signed(_GEN_539); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_541 = 5'h9 == _T_12 ? $signed(regsB_5_im) : $signed(_GEN_540); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_542 = 5'ha == _T_12 ? $signed(regsB_9_im) : $signed(_GEN_541); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_543 = 5'hb == _T_12 ? $signed(regsB_13_im) : $signed(_GEN_542); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_544 = 5'hc == _T_12 ? $signed(64'sh0) : $signed(_GEN_543); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_545 = 5'hd == _T_12 ? $signed(64'sh0) : $signed(_GEN_544); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_546 = 5'he == _T_12 ? $signed(64'sh0) : $signed(_GEN_545); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_547 = 5'hf == _T_12 ? $signed(64'sh0) : $signed(_GEN_546); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_548 = 5'h10 == _T_12 ? $signed(64'sh0) : $signed(_GEN_547); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_549 = 5'h11 == _T_12 ? $signed(64'sh0) : $signed(_GEN_548); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_550 = 5'h12 == _T_12 ? $signed(regsB_10_im) : $signed(_GEN_549); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_551 = 5'h13 == _T_12 ? $signed(regsB_14_im) : $signed(_GEN_550); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_552 = 5'h14 == _T_12 ? $signed(64'sh0) : $signed(_GEN_551); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_553 = 5'h15 == _T_12 ? $signed(64'sh0) : $signed(_GEN_552); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_554 = 5'h16 == _T_12 ? $signed(64'sh0) : $signed(_GEN_553); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_555 = 5'h17 == _T_12 ? $signed(64'sh0) : $signed(_GEN_554); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_556 = 5'h18 == _T_12 ? $signed(64'sh0) : $signed(_GEN_555); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_557 = 5'h19 == _T_12 ? $signed(64'sh0) : $signed(_GEN_556); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_558 = 5'h1a == _T_12 ? $signed(64'sh0) : $signed(_GEN_557); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_559 = 5'h1b == _T_12 ? $signed(regsB_15_im) : $signed(_GEN_558); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_561 = 5'h1 == _T_12 ? $signed(regsB_4_re) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_562 = 5'h2 == _T_12 ? $signed(regsB_8_re) : $signed(_GEN_561); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_563 = 5'h3 == _T_12 ? $signed(regsB_12_re) : $signed(_GEN_562); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_564 = 5'h4 == _T_12 ? $signed(64'sh0) : $signed(_GEN_563); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_565 = 5'h5 == _T_12 ? $signed(64'sh0) : $signed(_GEN_564); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_566 = 5'h6 == _T_12 ? $signed(64'sh0) : $signed(_GEN_565); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_567 = 5'h7 == _T_12 ? $signed(64'sh0) : $signed(_GEN_566); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_568 = 5'h8 == _T_12 ? $signed(64'sh0) : $signed(_GEN_567); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_569 = 5'h9 == _T_12 ? $signed(regsB_5_re) : $signed(_GEN_568); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_570 = 5'ha == _T_12 ? $signed(regsB_9_re) : $signed(_GEN_569); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_571 = 5'hb == _T_12 ? $signed(regsB_13_re) : $signed(_GEN_570); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_572 = 5'hc == _T_12 ? $signed(64'sh0) : $signed(_GEN_571); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_573 = 5'hd == _T_12 ? $signed(64'sh0) : $signed(_GEN_572); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_574 = 5'he == _T_12 ? $signed(64'sh0) : $signed(_GEN_573); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_575 = 5'hf == _T_12 ? $signed(64'sh0) : $signed(_GEN_574); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_576 = 5'h10 == _T_12 ? $signed(64'sh0) : $signed(_GEN_575); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_577 = 5'h11 == _T_12 ? $signed(64'sh0) : $signed(_GEN_576); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_578 = 5'h12 == _T_12 ? $signed(regsB_10_re) : $signed(_GEN_577); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_579 = 5'h13 == _T_12 ? $signed(regsB_14_re) : $signed(_GEN_578); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_580 = 5'h14 == _T_12 ? $signed(64'sh0) : $signed(_GEN_579); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_581 = 5'h15 == _T_12 ? $signed(64'sh0) : $signed(_GEN_580); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_582 = 5'h16 == _T_12 ? $signed(64'sh0) : $signed(_GEN_581); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_583 = 5'h17 == _T_12 ? $signed(64'sh0) : $signed(_GEN_582); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_584 = 5'h18 == _T_12 ? $signed(64'sh0) : $signed(_GEN_583); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_585 = 5'h19 == _T_12 ? $signed(64'sh0) : $signed(_GEN_584); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_586 = 5'h1a == _T_12 ? $signed(64'sh0) : $signed(_GEN_585); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_587 = 5'h1b == _T_12 ? $signed(regsB_15_re) : $signed(_GEN_586); // @[Matrix_Mul_V1.scala 162:{19,19}]
  PE PE ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_clock),
    .io_reset(PE_io_reset),
    .io_in_x_re(PE_io_in_x_re),
    .io_in_x_im(PE_io_in_x_im),
    .io_in_y_re(PE_io_in_y_re),
    .io_in_y_im(PE_io_in_y_im),
    .io_out_pe_re(PE_io_out_pe_re),
    .io_out_pe_im(PE_io_out_pe_im),
    .io_out_x_re(PE_io_out_x_re),
    .io_out_x_im(PE_io_out_x_im),
    .io_out_y_re(PE_io_out_y_re),
    .io_out_y_im(PE_io_out_y_im)
  );
  PE PE_1 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_1_clock),
    .io_reset(PE_1_io_reset),
    .io_in_x_re(PE_1_io_in_x_re),
    .io_in_x_im(PE_1_io_in_x_im),
    .io_in_y_re(PE_1_io_in_y_re),
    .io_in_y_im(PE_1_io_in_y_im),
    .io_out_pe_re(PE_1_io_out_pe_re),
    .io_out_pe_im(PE_1_io_out_pe_im),
    .io_out_x_re(PE_1_io_out_x_re),
    .io_out_x_im(PE_1_io_out_x_im),
    .io_out_y_re(PE_1_io_out_y_re),
    .io_out_y_im(PE_1_io_out_y_im)
  );
  PE PE_2 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_2_clock),
    .io_reset(PE_2_io_reset),
    .io_in_x_re(PE_2_io_in_x_re),
    .io_in_x_im(PE_2_io_in_x_im),
    .io_in_y_re(PE_2_io_in_y_re),
    .io_in_y_im(PE_2_io_in_y_im),
    .io_out_pe_re(PE_2_io_out_pe_re),
    .io_out_pe_im(PE_2_io_out_pe_im),
    .io_out_x_re(PE_2_io_out_x_re),
    .io_out_x_im(PE_2_io_out_x_im),
    .io_out_y_re(PE_2_io_out_y_re),
    .io_out_y_im(PE_2_io_out_y_im)
  );
  PE PE_3 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_3_clock),
    .io_reset(PE_3_io_reset),
    .io_in_x_re(PE_3_io_in_x_re),
    .io_in_x_im(PE_3_io_in_x_im),
    .io_in_y_re(PE_3_io_in_y_re),
    .io_in_y_im(PE_3_io_in_y_im),
    .io_out_pe_re(PE_3_io_out_pe_re),
    .io_out_pe_im(PE_3_io_out_pe_im),
    .io_out_x_re(PE_3_io_out_x_re),
    .io_out_x_im(PE_3_io_out_x_im),
    .io_out_y_re(PE_3_io_out_y_re),
    .io_out_y_im(PE_3_io_out_y_im)
  );
  PE PE_4 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_4_clock),
    .io_reset(PE_4_io_reset),
    .io_in_x_re(PE_4_io_in_x_re),
    .io_in_x_im(PE_4_io_in_x_im),
    .io_in_y_re(PE_4_io_in_y_re),
    .io_in_y_im(PE_4_io_in_y_im),
    .io_out_pe_re(PE_4_io_out_pe_re),
    .io_out_pe_im(PE_4_io_out_pe_im),
    .io_out_x_re(PE_4_io_out_x_re),
    .io_out_x_im(PE_4_io_out_x_im),
    .io_out_y_re(PE_4_io_out_y_re),
    .io_out_y_im(PE_4_io_out_y_im)
  );
  PE PE_5 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_5_clock),
    .io_reset(PE_5_io_reset),
    .io_in_x_re(PE_5_io_in_x_re),
    .io_in_x_im(PE_5_io_in_x_im),
    .io_in_y_re(PE_5_io_in_y_re),
    .io_in_y_im(PE_5_io_in_y_im),
    .io_out_pe_re(PE_5_io_out_pe_re),
    .io_out_pe_im(PE_5_io_out_pe_im),
    .io_out_x_re(PE_5_io_out_x_re),
    .io_out_x_im(PE_5_io_out_x_im),
    .io_out_y_re(PE_5_io_out_y_re),
    .io_out_y_im(PE_5_io_out_y_im)
  );
  PE PE_6 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_6_clock),
    .io_reset(PE_6_io_reset),
    .io_in_x_re(PE_6_io_in_x_re),
    .io_in_x_im(PE_6_io_in_x_im),
    .io_in_y_re(PE_6_io_in_y_re),
    .io_in_y_im(PE_6_io_in_y_im),
    .io_out_pe_re(PE_6_io_out_pe_re),
    .io_out_pe_im(PE_6_io_out_pe_im),
    .io_out_x_re(PE_6_io_out_x_re),
    .io_out_x_im(PE_6_io_out_x_im),
    .io_out_y_re(PE_6_io_out_y_re),
    .io_out_y_im(PE_6_io_out_y_im)
  );
  PE PE_7 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_7_clock),
    .io_reset(PE_7_io_reset),
    .io_in_x_re(PE_7_io_in_x_re),
    .io_in_x_im(PE_7_io_in_x_im),
    .io_in_y_re(PE_7_io_in_y_re),
    .io_in_y_im(PE_7_io_in_y_im),
    .io_out_pe_re(PE_7_io_out_pe_re),
    .io_out_pe_im(PE_7_io_out_pe_im),
    .io_out_x_re(PE_7_io_out_x_re),
    .io_out_x_im(PE_7_io_out_x_im),
    .io_out_y_re(PE_7_io_out_y_re),
    .io_out_y_im(PE_7_io_out_y_im)
  );
  PE PE_8 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_8_clock),
    .io_reset(PE_8_io_reset),
    .io_in_x_re(PE_8_io_in_x_re),
    .io_in_x_im(PE_8_io_in_x_im),
    .io_in_y_re(PE_8_io_in_y_re),
    .io_in_y_im(PE_8_io_in_y_im),
    .io_out_pe_re(PE_8_io_out_pe_re),
    .io_out_pe_im(PE_8_io_out_pe_im),
    .io_out_x_re(PE_8_io_out_x_re),
    .io_out_x_im(PE_8_io_out_x_im),
    .io_out_y_re(PE_8_io_out_y_re),
    .io_out_y_im(PE_8_io_out_y_im)
  );
  PE PE_9 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_9_clock),
    .io_reset(PE_9_io_reset),
    .io_in_x_re(PE_9_io_in_x_re),
    .io_in_x_im(PE_9_io_in_x_im),
    .io_in_y_re(PE_9_io_in_y_re),
    .io_in_y_im(PE_9_io_in_y_im),
    .io_out_pe_re(PE_9_io_out_pe_re),
    .io_out_pe_im(PE_9_io_out_pe_im),
    .io_out_x_re(PE_9_io_out_x_re),
    .io_out_x_im(PE_9_io_out_x_im),
    .io_out_y_re(PE_9_io_out_y_re),
    .io_out_y_im(PE_9_io_out_y_im)
  );
  PE PE_10 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_10_clock),
    .io_reset(PE_10_io_reset),
    .io_in_x_re(PE_10_io_in_x_re),
    .io_in_x_im(PE_10_io_in_x_im),
    .io_in_y_re(PE_10_io_in_y_re),
    .io_in_y_im(PE_10_io_in_y_im),
    .io_out_pe_re(PE_10_io_out_pe_re),
    .io_out_pe_im(PE_10_io_out_pe_im),
    .io_out_x_re(PE_10_io_out_x_re),
    .io_out_x_im(PE_10_io_out_x_im),
    .io_out_y_re(PE_10_io_out_y_re),
    .io_out_y_im(PE_10_io_out_y_im)
  );
  PE PE_11 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_11_clock),
    .io_reset(PE_11_io_reset),
    .io_in_x_re(PE_11_io_in_x_re),
    .io_in_x_im(PE_11_io_in_x_im),
    .io_in_y_re(PE_11_io_in_y_re),
    .io_in_y_im(PE_11_io_in_y_im),
    .io_out_pe_re(PE_11_io_out_pe_re),
    .io_out_pe_im(PE_11_io_out_pe_im),
    .io_out_x_re(PE_11_io_out_x_re),
    .io_out_x_im(PE_11_io_out_x_im),
    .io_out_y_re(PE_11_io_out_y_re),
    .io_out_y_im(PE_11_io_out_y_im)
  );
  PE PE_12 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_12_clock),
    .io_reset(PE_12_io_reset),
    .io_in_x_re(PE_12_io_in_x_re),
    .io_in_x_im(PE_12_io_in_x_im),
    .io_in_y_re(PE_12_io_in_y_re),
    .io_in_y_im(PE_12_io_in_y_im),
    .io_out_pe_re(PE_12_io_out_pe_re),
    .io_out_pe_im(PE_12_io_out_pe_im),
    .io_out_x_re(PE_12_io_out_x_re),
    .io_out_x_im(PE_12_io_out_x_im),
    .io_out_y_re(PE_12_io_out_y_re),
    .io_out_y_im(PE_12_io_out_y_im)
  );
  PE PE_13 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_13_clock),
    .io_reset(PE_13_io_reset),
    .io_in_x_re(PE_13_io_in_x_re),
    .io_in_x_im(PE_13_io_in_x_im),
    .io_in_y_re(PE_13_io_in_y_re),
    .io_in_y_im(PE_13_io_in_y_im),
    .io_out_pe_re(PE_13_io_out_pe_re),
    .io_out_pe_im(PE_13_io_out_pe_im),
    .io_out_x_re(PE_13_io_out_x_re),
    .io_out_x_im(PE_13_io_out_x_im),
    .io_out_y_re(PE_13_io_out_y_re),
    .io_out_y_im(PE_13_io_out_y_im)
  );
  PE PE_14 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_14_clock),
    .io_reset(PE_14_io_reset),
    .io_in_x_re(PE_14_io_in_x_re),
    .io_in_x_im(PE_14_io_in_x_im),
    .io_in_y_re(PE_14_io_in_y_re),
    .io_in_y_im(PE_14_io_in_y_im),
    .io_out_pe_re(PE_14_io_out_pe_re),
    .io_out_pe_im(PE_14_io_out_pe_im),
    .io_out_x_re(PE_14_io_out_x_re),
    .io_out_x_im(PE_14_io_out_x_im),
    .io_out_y_re(PE_14_io_out_y_re),
    .io_out_y_im(PE_14_io_out_y_im)
  );
  PE PE_15 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_15_clock),
    .io_reset(PE_15_io_reset),
    .io_in_x_re(PE_15_io_in_x_re),
    .io_in_x_im(PE_15_io_in_x_im),
    .io_in_y_re(PE_15_io_in_y_re),
    .io_in_y_im(PE_15_io_in_y_im),
    .io_out_pe_re(PE_15_io_out_pe_re),
    .io_out_pe_im(PE_15_io_out_pe_im),
    .io_out_x_re(PE_15_io_out_x_re),
    .io_out_x_im(PE_15_io_out_x_im),
    .io_out_y_re(PE_15_io_out_y_re),
    .io_out_y_im(PE_15_io_out_y_im)
  );
  assign io_matrixC_0_re = PE_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_0_im = PE_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_1_re = PE_1_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_1_im = PE_1_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_2_re = PE_2_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_2_im = PE_2_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_3_re = PE_3_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_3_im = PE_3_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_4_re = PE_4_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_4_im = PE_4_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_5_re = PE_5_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_5_im = PE_5_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_6_re = PE_6_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_6_im = PE_6_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_7_re = PE_7_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_7_im = PE_7_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_8_re = PE_8_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_8_im = PE_8_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_9_re = PE_9_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_9_im = PE_9_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_10_re = PE_10_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_10_im = PE_10_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_11_re = PE_11_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_11_im = PE_11_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_12_re = PE_12_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_12_im = PE_12_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_13_re = PE_13_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_13_im = PE_13_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_14_re = PE_14_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_14_im = PE_14_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_15_re = PE_15_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_15_im = PE_15_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_valid = input_point >= 5'ha; // @[Matrix_Mul_V1.scala 188:20]
  assign PE_clock = clock;
  assign PE_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_io_in_x_re = input_point < 5'h7 ? $signed(_GEN_187) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_io_in_x_im = input_point < 5'h7 ? $signed(_GEN_159) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_io_in_y_re = _T ? $signed(_GEN_419) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_io_in_y_im = _T ? $signed(_GEN_391) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_1_clock = clock;
  assign PE_1_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_1_io_in_x_re = PE_io_out_x_re; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_1_io_in_x_im = PE_io_out_x_im; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_1_io_in_y_re = _T ? $signed(_GEN_475) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_1_io_in_y_im = _T ? $signed(_GEN_447) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_2_clock = clock;
  assign PE_2_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_2_io_in_x_re = PE_1_io_out_x_re; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_2_io_in_x_im = PE_1_io_out_x_im; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_2_io_in_y_re = _T ? $signed(_GEN_531) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_2_io_in_y_im = _T ? $signed(_GEN_503) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_3_clock = clock;
  assign PE_3_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_3_io_in_x_re = PE_2_io_out_x_re; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_3_io_in_x_im = PE_2_io_out_x_im; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_3_io_in_y_re = _T ? $signed(_GEN_587) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_3_io_in_y_im = _T ? $signed(_GEN_559) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_4_clock = clock;
  assign PE_4_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_4_io_in_x_re = input_point < 5'h7 ? $signed(_GEN_243) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_4_io_in_x_im = input_point < 5'h7 ? $signed(_GEN_215) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_4_io_in_y_re = PE_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_4_io_in_y_im = PE_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_5_clock = clock;
  assign PE_5_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_5_io_in_x_re = PE_4_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_5_io_in_x_im = PE_4_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_5_io_in_y_re = PE_1_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_5_io_in_y_im = PE_1_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_6_clock = clock;
  assign PE_6_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_6_io_in_x_re = PE_5_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_6_io_in_x_im = PE_5_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_6_io_in_y_re = PE_2_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_6_io_in_y_im = PE_2_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_7_clock = clock;
  assign PE_7_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_7_io_in_x_re = PE_6_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_7_io_in_x_im = PE_6_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_7_io_in_y_re = PE_3_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_7_io_in_y_im = PE_3_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_8_clock = clock;
  assign PE_8_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_8_io_in_x_re = input_point < 5'h7 ? $signed(_GEN_299) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_8_io_in_x_im = input_point < 5'h7 ? $signed(_GEN_271) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_8_io_in_y_re = PE_4_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_8_io_in_y_im = PE_4_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_9_clock = clock;
  assign PE_9_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_9_io_in_x_re = PE_8_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_9_io_in_x_im = PE_8_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_9_io_in_y_re = PE_5_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_9_io_in_y_im = PE_5_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_10_clock = clock;
  assign PE_10_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_10_io_in_x_re = PE_9_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_10_io_in_x_im = PE_9_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_10_io_in_y_re = PE_6_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_10_io_in_y_im = PE_6_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_11_clock = clock;
  assign PE_11_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_11_io_in_x_re = PE_10_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_11_io_in_x_im = PE_10_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_11_io_in_y_re = PE_7_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_11_io_in_y_im = PE_7_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_12_clock = clock;
  assign PE_12_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_12_io_in_x_re = input_point < 5'h7 ? $signed(_GEN_355) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_12_io_in_x_im = input_point < 5'h7 ? $signed(_GEN_327) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_12_io_in_y_re = PE_8_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_12_io_in_y_im = PE_8_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_13_clock = clock;
  assign PE_13_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_13_io_in_x_re = PE_12_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_13_io_in_x_im = PE_12_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_13_io_in_y_re = PE_9_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_13_io_in_y_im = PE_9_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_14_clock = clock;
  assign PE_14_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_14_io_in_x_re = PE_13_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_14_io_in_x_im = PE_13_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_14_io_in_y_re = PE_10_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_14_io_in_y_im = PE_10_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_15_clock = clock;
  assign PE_15_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_15_io_in_x_re = PE_14_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_15_io_in_x_im = PE_14_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_15_io_in_y_re = PE_11_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_15_io_in_y_im = PE_11_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  always @(posedge clock) begin
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_0_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_0_re <= io_matrixA_0_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_0_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_0_im <= io_matrixA_0_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_1_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_1_re <= io_matrixA_1_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_1_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_1_im <= io_matrixA_1_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_2_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_2_re <= io_matrixA_2_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_2_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_2_im <= io_matrixA_2_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_3_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_3_re <= io_matrixA_3_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_3_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_3_im <= io_matrixA_3_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_5_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_5_re <= io_matrixA_5_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_5_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_5_im <= io_matrixA_5_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_6_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_6_re <= io_matrixA_6_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_6_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_6_im <= io_matrixA_6_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_7_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_7_re <= io_matrixA_7_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_7_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_7_im <= io_matrixA_7_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_10_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_10_re <= io_matrixA_10_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_10_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_10_im <= io_matrixA_10_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_11_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_11_re <= io_matrixA_11_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_11_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_11_im <= io_matrixA_11_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_15_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_15_re <= io_matrixA_15_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_15_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_15_im <= io_matrixA_15_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_0_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_0_re <= io_matrixB_0_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_0_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_0_im <= io_matrixB_0_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_4_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_4_re <= io_matrixB_4_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_4_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_4_im <= io_matrixB_4_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_5_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_5_re <= io_matrixB_5_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_5_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_5_im <= io_matrixB_5_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_8_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_8_re <= io_matrixB_8_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_8_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_8_im <= io_matrixB_8_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_9_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_9_re <= io_matrixB_9_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_9_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_9_im <= io_matrixB_9_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_10_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_10_re <= io_matrixB_10_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_10_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_10_im <= io_matrixB_10_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_12_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_12_re <= io_matrixB_12_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_12_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_12_im <= io_matrixB_12_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_13_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_13_re <= io_matrixB_13_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_13_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_13_im <= io_matrixB_13_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_14_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_14_re <= io_matrixB_14_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_14_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_14_im <= io_matrixB_14_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_15_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_15_re <= io_matrixB_15_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_15_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_15_im <= io_matrixB_15_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      input_point <= 5'h0; // @[Matrix_Mul_V1.scala 99:17]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      input_point <= 5'h0; // @[Matrix_Mul_V1.scala 108:17]
    end else begin
      input_point <= _input_point_T_1; // @[Matrix_Mul_V1.scala 116:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regsA_0_re = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regsA_0_im = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  regsA_1_re = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  regsA_1_im = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  regsA_2_re = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  regsA_2_im = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  regsA_3_re = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  regsA_3_im = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  regsA_5_re = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  regsA_5_im = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  regsA_6_re = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  regsA_6_im = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  regsA_7_re = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  regsA_7_im = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  regsA_10_re = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  regsA_10_im = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  regsA_11_re = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  regsA_11_im = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  regsA_15_re = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  regsA_15_im = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  regsB_0_re = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  regsB_0_im = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  regsB_4_re = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  regsB_4_im = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  regsB_5_re = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  regsB_5_im = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  regsB_8_re = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  regsB_8_im = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  regsB_9_re = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  regsB_9_im = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  regsB_10_re = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  regsB_10_im = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  regsB_12_re = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  regsB_12_im = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  regsB_13_re = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  regsB_13_im = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  regsB_14_re = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  regsB_14_im = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  regsB_15_re = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  regsB_15_im = _RAND_39[63:0];
  _RAND_40 = {1{`RANDOM}};
  input_point = _RAND_40[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module matrix_mul_v1_3(
  input         clock,
  input         io_reset,
  input         io_ready,
  input  [63:0] io_matrixA_0_re,
  input  [63:0] io_matrixA_0_im,
  input  [63:0] io_matrixA_1_re,
  input  [63:0] io_matrixA_1_im,
  input  [63:0] io_matrixA_2_re,
  input  [63:0] io_matrixA_2_im,
  input  [63:0] io_matrixA_3_re,
  input  [63:0] io_matrixA_3_im,
  input  [63:0] io_matrixA_4_re,
  input  [63:0] io_matrixA_4_im,
  input  [63:0] io_matrixA_5_re,
  input  [63:0] io_matrixA_5_im,
  input  [63:0] io_matrixA_6_re,
  input  [63:0] io_matrixA_6_im,
  input  [63:0] io_matrixA_7_re,
  input  [63:0] io_matrixA_7_im,
  input  [63:0] io_matrixA_8_re,
  input  [63:0] io_matrixA_8_im,
  input  [63:0] io_matrixA_9_re,
  input  [63:0] io_matrixA_9_im,
  input  [63:0] io_matrixA_10_re,
  input  [63:0] io_matrixA_10_im,
  input  [63:0] io_matrixA_11_re,
  input  [63:0] io_matrixA_11_im,
  input  [63:0] io_matrixA_12_re,
  input  [63:0] io_matrixA_12_im,
  input  [63:0] io_matrixA_13_re,
  input  [63:0] io_matrixA_13_im,
  input  [63:0] io_matrixA_14_re,
  input  [63:0] io_matrixA_14_im,
  input  [63:0] io_matrixA_15_re,
  input  [63:0] io_matrixA_15_im,
  input  [63:0] io_matrixB_0_re,
  input  [63:0] io_matrixB_0_im,
  input  [63:0] io_matrixB_1_re,
  input  [63:0] io_matrixB_1_im,
  input  [63:0] io_matrixB_2_re,
  input  [63:0] io_matrixB_2_im,
  input  [63:0] io_matrixB_3_re,
  input  [63:0] io_matrixB_3_im,
  output [63:0] io_matrixC_0_re,
  output [63:0] io_matrixC_0_im,
  output [63:0] io_matrixC_1_re,
  output [63:0] io_matrixC_1_im,
  output [63:0] io_matrixC_2_re,
  output [63:0] io_matrixC_2_im,
  output [63:0] io_matrixC_3_re,
  output [63:0] io_matrixC_3_im,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [31:0] _RAND_40;
`endif // RANDOMIZE_REG_INIT
  wire  PE_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_1_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_1_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_1_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_2_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_2_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_2_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_3_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_3_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [63:0] PE_3_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  reg [63:0] regsA_0_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_0_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_1_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_1_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_2_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_2_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_3_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_3_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_4_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_4_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_5_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_5_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_6_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_6_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_7_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_7_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_8_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_8_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_9_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_9_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_10_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_10_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_11_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_11_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_12_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_12_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_13_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_13_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_14_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_14_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_15_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsA_15_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [63:0] regsB_0_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_0_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_1_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_1_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_2_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_2_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_3_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [63:0] regsB_3_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [4:0] input_point; // @[Matrix_Mul_V1.scala 84:30]
  wire [4:0] _input_point_T_1 = input_point + 5'h1; // @[Matrix_Mul_V1.scala 116:32]
  wire [3:0] _T_1 = 1'h0 * 3'h7; // @[Matrix_Mul_V1.scala 148:44]
  wire [4:0] _GEN_327 = {{1'd0}, _T_1}; // @[Matrix_Mul_V1.scala 148:60]
  wire [4:0] _T_3 = _GEN_327 + input_point; // @[Matrix_Mul_V1.scala 148:60]
  wire [63:0] _GEN_85 = 5'h1 == _T_3 ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_86 = 5'h2 == _T_3 ? $signed(regsA_2_im) : $signed(_GEN_85); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_87 = 5'h3 == _T_3 ? $signed(regsA_3_im) : $signed(_GEN_86); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_88 = 5'h4 == _T_3 ? $signed(64'sh0) : $signed(_GEN_87); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_89 = 5'h5 == _T_3 ? $signed(64'sh0) : $signed(_GEN_88); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_90 = 5'h6 == _T_3 ? $signed(64'sh0) : $signed(_GEN_89); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_91 = 5'h7 == _T_3 ? $signed(64'sh0) : $signed(_GEN_90); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_92 = 5'h8 == _T_3 ? $signed(regsA_4_im) : $signed(_GEN_91); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_93 = 5'h9 == _T_3 ? $signed(regsA_5_im) : $signed(_GEN_92); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_94 = 5'ha == _T_3 ? $signed(regsA_6_im) : $signed(_GEN_93); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_95 = 5'hb == _T_3 ? $signed(regsA_7_im) : $signed(_GEN_94); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_96 = 5'hc == _T_3 ? $signed(64'sh0) : $signed(_GEN_95); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_97 = 5'hd == _T_3 ? $signed(64'sh0) : $signed(_GEN_96); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_98 = 5'he == _T_3 ? $signed(64'sh0) : $signed(_GEN_97); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_99 = 5'hf == _T_3 ? $signed(64'sh0) : $signed(_GEN_98); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_100 = 5'h10 == _T_3 ? $signed(regsA_8_im) : $signed(_GEN_99); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_101 = 5'h11 == _T_3 ? $signed(regsA_9_im) : $signed(_GEN_100); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_102 = 5'h12 == _T_3 ? $signed(regsA_10_im) : $signed(_GEN_101); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_103 = 5'h13 == _T_3 ? $signed(regsA_11_im) : $signed(_GEN_102); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_104 = 5'h14 == _T_3 ? $signed(64'sh0) : $signed(_GEN_103); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_105 = 5'h15 == _T_3 ? $signed(64'sh0) : $signed(_GEN_104); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_106 = 5'h16 == _T_3 ? $signed(64'sh0) : $signed(_GEN_105); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_107 = 5'h17 == _T_3 ? $signed(64'sh0) : $signed(_GEN_106); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_108 = 5'h18 == _T_3 ? $signed(regsA_12_im) : $signed(_GEN_107); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_109 = 5'h19 == _T_3 ? $signed(regsA_13_im) : $signed(_GEN_108); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_110 = 5'h1a == _T_3 ? $signed(regsA_14_im) : $signed(_GEN_109); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_111 = 5'h1b == _T_3 ? $signed(regsA_15_im) : $signed(_GEN_110); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_113 = 5'h1 == _T_3 ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_114 = 5'h2 == _T_3 ? $signed(regsA_2_re) : $signed(_GEN_113); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_115 = 5'h3 == _T_3 ? $signed(regsA_3_re) : $signed(_GEN_114); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_116 = 5'h4 == _T_3 ? $signed(64'sh0) : $signed(_GEN_115); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_117 = 5'h5 == _T_3 ? $signed(64'sh0) : $signed(_GEN_116); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_118 = 5'h6 == _T_3 ? $signed(64'sh0) : $signed(_GEN_117); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_119 = 5'h7 == _T_3 ? $signed(64'sh0) : $signed(_GEN_118); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_120 = 5'h8 == _T_3 ? $signed(regsA_4_re) : $signed(_GEN_119); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_121 = 5'h9 == _T_3 ? $signed(regsA_5_re) : $signed(_GEN_120); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_122 = 5'ha == _T_3 ? $signed(regsA_6_re) : $signed(_GEN_121); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_123 = 5'hb == _T_3 ? $signed(regsA_7_re) : $signed(_GEN_122); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_124 = 5'hc == _T_3 ? $signed(64'sh0) : $signed(_GEN_123); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_125 = 5'hd == _T_3 ? $signed(64'sh0) : $signed(_GEN_124); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_126 = 5'he == _T_3 ? $signed(64'sh0) : $signed(_GEN_125); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_127 = 5'hf == _T_3 ? $signed(64'sh0) : $signed(_GEN_126); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_128 = 5'h10 == _T_3 ? $signed(regsA_8_re) : $signed(_GEN_127); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_129 = 5'h11 == _T_3 ? $signed(regsA_9_re) : $signed(_GEN_128); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_130 = 5'h12 == _T_3 ? $signed(regsA_10_re) : $signed(_GEN_129); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_131 = 5'h13 == _T_3 ? $signed(regsA_11_re) : $signed(_GEN_130); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_132 = 5'h14 == _T_3 ? $signed(64'sh0) : $signed(_GEN_131); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_133 = 5'h15 == _T_3 ? $signed(64'sh0) : $signed(_GEN_132); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_134 = 5'h16 == _T_3 ? $signed(64'sh0) : $signed(_GEN_133); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_135 = 5'h17 == _T_3 ? $signed(64'sh0) : $signed(_GEN_134); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_136 = 5'h18 == _T_3 ? $signed(regsA_12_re) : $signed(_GEN_135); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_137 = 5'h19 == _T_3 ? $signed(regsA_13_re) : $signed(_GEN_136); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_138 = 5'h1a == _T_3 ? $signed(regsA_14_re) : $signed(_GEN_137); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_139 = 5'h1b == _T_3 ? $signed(regsA_15_re) : $signed(_GEN_138); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [3:0] _T_4 = 1'h1 * 3'h7; // @[Matrix_Mul_V1.scala 148:44]
  wire [4:0] _GEN_328 = {{1'd0}, _T_4}; // @[Matrix_Mul_V1.scala 148:60]
  wire [4:0] _T_6 = _GEN_328 + input_point; // @[Matrix_Mul_V1.scala 148:60]
  wire [63:0] _GEN_141 = 5'h1 == _T_6 ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_142 = 5'h2 == _T_6 ? $signed(regsA_2_im) : $signed(_GEN_141); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_143 = 5'h3 == _T_6 ? $signed(regsA_3_im) : $signed(_GEN_142); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_144 = 5'h4 == _T_6 ? $signed(64'sh0) : $signed(_GEN_143); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_145 = 5'h5 == _T_6 ? $signed(64'sh0) : $signed(_GEN_144); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_146 = 5'h6 == _T_6 ? $signed(64'sh0) : $signed(_GEN_145); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_147 = 5'h7 == _T_6 ? $signed(64'sh0) : $signed(_GEN_146); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_148 = 5'h8 == _T_6 ? $signed(regsA_4_im) : $signed(_GEN_147); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_149 = 5'h9 == _T_6 ? $signed(regsA_5_im) : $signed(_GEN_148); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_150 = 5'ha == _T_6 ? $signed(regsA_6_im) : $signed(_GEN_149); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_151 = 5'hb == _T_6 ? $signed(regsA_7_im) : $signed(_GEN_150); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_152 = 5'hc == _T_6 ? $signed(64'sh0) : $signed(_GEN_151); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_153 = 5'hd == _T_6 ? $signed(64'sh0) : $signed(_GEN_152); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_154 = 5'he == _T_6 ? $signed(64'sh0) : $signed(_GEN_153); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_155 = 5'hf == _T_6 ? $signed(64'sh0) : $signed(_GEN_154); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_156 = 5'h10 == _T_6 ? $signed(regsA_8_im) : $signed(_GEN_155); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_157 = 5'h11 == _T_6 ? $signed(regsA_9_im) : $signed(_GEN_156); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_158 = 5'h12 == _T_6 ? $signed(regsA_10_im) : $signed(_GEN_157); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_159 = 5'h13 == _T_6 ? $signed(regsA_11_im) : $signed(_GEN_158); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_160 = 5'h14 == _T_6 ? $signed(64'sh0) : $signed(_GEN_159); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_161 = 5'h15 == _T_6 ? $signed(64'sh0) : $signed(_GEN_160); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_162 = 5'h16 == _T_6 ? $signed(64'sh0) : $signed(_GEN_161); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_163 = 5'h17 == _T_6 ? $signed(64'sh0) : $signed(_GEN_162); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_164 = 5'h18 == _T_6 ? $signed(regsA_12_im) : $signed(_GEN_163); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_165 = 5'h19 == _T_6 ? $signed(regsA_13_im) : $signed(_GEN_164); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_166 = 5'h1a == _T_6 ? $signed(regsA_14_im) : $signed(_GEN_165); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_167 = 5'h1b == _T_6 ? $signed(regsA_15_im) : $signed(_GEN_166); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_169 = 5'h1 == _T_6 ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_170 = 5'h2 == _T_6 ? $signed(regsA_2_re) : $signed(_GEN_169); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_171 = 5'h3 == _T_6 ? $signed(regsA_3_re) : $signed(_GEN_170); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_172 = 5'h4 == _T_6 ? $signed(64'sh0) : $signed(_GEN_171); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_173 = 5'h5 == _T_6 ? $signed(64'sh0) : $signed(_GEN_172); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_174 = 5'h6 == _T_6 ? $signed(64'sh0) : $signed(_GEN_173); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_175 = 5'h7 == _T_6 ? $signed(64'sh0) : $signed(_GEN_174); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_176 = 5'h8 == _T_6 ? $signed(regsA_4_re) : $signed(_GEN_175); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_177 = 5'h9 == _T_6 ? $signed(regsA_5_re) : $signed(_GEN_176); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_178 = 5'ha == _T_6 ? $signed(regsA_6_re) : $signed(_GEN_177); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_179 = 5'hb == _T_6 ? $signed(regsA_7_re) : $signed(_GEN_178); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_180 = 5'hc == _T_6 ? $signed(64'sh0) : $signed(_GEN_179); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_181 = 5'hd == _T_6 ? $signed(64'sh0) : $signed(_GEN_180); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_182 = 5'he == _T_6 ? $signed(64'sh0) : $signed(_GEN_181); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_183 = 5'hf == _T_6 ? $signed(64'sh0) : $signed(_GEN_182); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_184 = 5'h10 == _T_6 ? $signed(regsA_8_re) : $signed(_GEN_183); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_185 = 5'h11 == _T_6 ? $signed(regsA_9_re) : $signed(_GEN_184); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_186 = 5'h12 == _T_6 ? $signed(regsA_10_re) : $signed(_GEN_185); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_187 = 5'h13 == _T_6 ? $signed(regsA_11_re) : $signed(_GEN_186); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_188 = 5'h14 == _T_6 ? $signed(64'sh0) : $signed(_GEN_187); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_189 = 5'h15 == _T_6 ? $signed(64'sh0) : $signed(_GEN_188); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_190 = 5'h16 == _T_6 ? $signed(64'sh0) : $signed(_GEN_189); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_191 = 5'h17 == _T_6 ? $signed(64'sh0) : $signed(_GEN_190); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_192 = 5'h18 == _T_6 ? $signed(regsA_12_re) : $signed(_GEN_191); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_193 = 5'h19 == _T_6 ? $signed(regsA_13_re) : $signed(_GEN_192); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_194 = 5'h1a == _T_6 ? $signed(regsA_14_re) : $signed(_GEN_193); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_195 = 5'h1b == _T_6 ? $signed(regsA_15_re) : $signed(_GEN_194); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [4:0] _T_7 = 2'h2 * 3'h7; // @[Matrix_Mul_V1.scala 148:44]
  wire [4:0] _T_9 = _T_7 + input_point; // @[Matrix_Mul_V1.scala 148:60]
  wire [63:0] _GEN_197 = 5'h1 == _T_9 ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_198 = 5'h2 == _T_9 ? $signed(regsA_2_im) : $signed(_GEN_197); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_199 = 5'h3 == _T_9 ? $signed(regsA_3_im) : $signed(_GEN_198); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_200 = 5'h4 == _T_9 ? $signed(64'sh0) : $signed(_GEN_199); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_201 = 5'h5 == _T_9 ? $signed(64'sh0) : $signed(_GEN_200); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_202 = 5'h6 == _T_9 ? $signed(64'sh0) : $signed(_GEN_201); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_203 = 5'h7 == _T_9 ? $signed(64'sh0) : $signed(_GEN_202); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_204 = 5'h8 == _T_9 ? $signed(regsA_4_im) : $signed(_GEN_203); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_205 = 5'h9 == _T_9 ? $signed(regsA_5_im) : $signed(_GEN_204); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_206 = 5'ha == _T_9 ? $signed(regsA_6_im) : $signed(_GEN_205); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_207 = 5'hb == _T_9 ? $signed(regsA_7_im) : $signed(_GEN_206); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_208 = 5'hc == _T_9 ? $signed(64'sh0) : $signed(_GEN_207); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_209 = 5'hd == _T_9 ? $signed(64'sh0) : $signed(_GEN_208); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_210 = 5'he == _T_9 ? $signed(64'sh0) : $signed(_GEN_209); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_211 = 5'hf == _T_9 ? $signed(64'sh0) : $signed(_GEN_210); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_212 = 5'h10 == _T_9 ? $signed(regsA_8_im) : $signed(_GEN_211); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_213 = 5'h11 == _T_9 ? $signed(regsA_9_im) : $signed(_GEN_212); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_214 = 5'h12 == _T_9 ? $signed(regsA_10_im) : $signed(_GEN_213); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_215 = 5'h13 == _T_9 ? $signed(regsA_11_im) : $signed(_GEN_214); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_216 = 5'h14 == _T_9 ? $signed(64'sh0) : $signed(_GEN_215); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_217 = 5'h15 == _T_9 ? $signed(64'sh0) : $signed(_GEN_216); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_218 = 5'h16 == _T_9 ? $signed(64'sh0) : $signed(_GEN_217); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_219 = 5'h17 == _T_9 ? $signed(64'sh0) : $signed(_GEN_218); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_220 = 5'h18 == _T_9 ? $signed(regsA_12_im) : $signed(_GEN_219); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_221 = 5'h19 == _T_9 ? $signed(regsA_13_im) : $signed(_GEN_220); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_222 = 5'h1a == _T_9 ? $signed(regsA_14_im) : $signed(_GEN_221); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_223 = 5'h1b == _T_9 ? $signed(regsA_15_im) : $signed(_GEN_222); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_225 = 5'h1 == _T_9 ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_226 = 5'h2 == _T_9 ? $signed(regsA_2_re) : $signed(_GEN_225); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_227 = 5'h3 == _T_9 ? $signed(regsA_3_re) : $signed(_GEN_226); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_228 = 5'h4 == _T_9 ? $signed(64'sh0) : $signed(_GEN_227); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_229 = 5'h5 == _T_9 ? $signed(64'sh0) : $signed(_GEN_228); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_230 = 5'h6 == _T_9 ? $signed(64'sh0) : $signed(_GEN_229); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_231 = 5'h7 == _T_9 ? $signed(64'sh0) : $signed(_GEN_230); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_232 = 5'h8 == _T_9 ? $signed(regsA_4_re) : $signed(_GEN_231); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_233 = 5'h9 == _T_9 ? $signed(regsA_5_re) : $signed(_GEN_232); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_234 = 5'ha == _T_9 ? $signed(regsA_6_re) : $signed(_GEN_233); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_235 = 5'hb == _T_9 ? $signed(regsA_7_re) : $signed(_GEN_234); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_236 = 5'hc == _T_9 ? $signed(64'sh0) : $signed(_GEN_235); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_237 = 5'hd == _T_9 ? $signed(64'sh0) : $signed(_GEN_236); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_238 = 5'he == _T_9 ? $signed(64'sh0) : $signed(_GEN_237); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_239 = 5'hf == _T_9 ? $signed(64'sh0) : $signed(_GEN_238); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_240 = 5'h10 == _T_9 ? $signed(regsA_8_re) : $signed(_GEN_239); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_241 = 5'h11 == _T_9 ? $signed(regsA_9_re) : $signed(_GEN_240); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_242 = 5'h12 == _T_9 ? $signed(regsA_10_re) : $signed(_GEN_241); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_243 = 5'h13 == _T_9 ? $signed(regsA_11_re) : $signed(_GEN_242); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_244 = 5'h14 == _T_9 ? $signed(64'sh0) : $signed(_GEN_243); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_245 = 5'h15 == _T_9 ? $signed(64'sh0) : $signed(_GEN_244); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_246 = 5'h16 == _T_9 ? $signed(64'sh0) : $signed(_GEN_245); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_247 = 5'h17 == _T_9 ? $signed(64'sh0) : $signed(_GEN_246); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_248 = 5'h18 == _T_9 ? $signed(regsA_12_re) : $signed(_GEN_247); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_249 = 5'h19 == _T_9 ? $signed(regsA_13_re) : $signed(_GEN_248); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_250 = 5'h1a == _T_9 ? $signed(regsA_14_re) : $signed(_GEN_249); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_251 = 5'h1b == _T_9 ? $signed(regsA_15_re) : $signed(_GEN_250); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [4:0] _T_10 = 2'h3 * 3'h7; // @[Matrix_Mul_V1.scala 148:44]
  wire [4:0] _T_12 = _T_10 + input_point; // @[Matrix_Mul_V1.scala 148:60]
  wire [63:0] _GEN_253 = 5'h1 == _T_12 ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_254 = 5'h2 == _T_12 ? $signed(regsA_2_im) : $signed(_GEN_253); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_255 = 5'h3 == _T_12 ? $signed(regsA_3_im) : $signed(_GEN_254); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_256 = 5'h4 == _T_12 ? $signed(64'sh0) : $signed(_GEN_255); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_257 = 5'h5 == _T_12 ? $signed(64'sh0) : $signed(_GEN_256); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_258 = 5'h6 == _T_12 ? $signed(64'sh0) : $signed(_GEN_257); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_259 = 5'h7 == _T_12 ? $signed(64'sh0) : $signed(_GEN_258); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_260 = 5'h8 == _T_12 ? $signed(regsA_4_im) : $signed(_GEN_259); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_261 = 5'h9 == _T_12 ? $signed(regsA_5_im) : $signed(_GEN_260); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_262 = 5'ha == _T_12 ? $signed(regsA_6_im) : $signed(_GEN_261); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_263 = 5'hb == _T_12 ? $signed(regsA_7_im) : $signed(_GEN_262); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_264 = 5'hc == _T_12 ? $signed(64'sh0) : $signed(_GEN_263); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_265 = 5'hd == _T_12 ? $signed(64'sh0) : $signed(_GEN_264); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_266 = 5'he == _T_12 ? $signed(64'sh0) : $signed(_GEN_265); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_267 = 5'hf == _T_12 ? $signed(64'sh0) : $signed(_GEN_266); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_268 = 5'h10 == _T_12 ? $signed(regsA_8_im) : $signed(_GEN_267); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_269 = 5'h11 == _T_12 ? $signed(regsA_9_im) : $signed(_GEN_268); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_270 = 5'h12 == _T_12 ? $signed(regsA_10_im) : $signed(_GEN_269); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_271 = 5'h13 == _T_12 ? $signed(regsA_11_im) : $signed(_GEN_270); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_272 = 5'h14 == _T_12 ? $signed(64'sh0) : $signed(_GEN_271); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_273 = 5'h15 == _T_12 ? $signed(64'sh0) : $signed(_GEN_272); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_274 = 5'h16 == _T_12 ? $signed(64'sh0) : $signed(_GEN_273); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_275 = 5'h17 == _T_12 ? $signed(64'sh0) : $signed(_GEN_274); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_276 = 5'h18 == _T_12 ? $signed(regsA_12_im) : $signed(_GEN_275); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_277 = 5'h19 == _T_12 ? $signed(regsA_13_im) : $signed(_GEN_276); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_278 = 5'h1a == _T_12 ? $signed(regsA_14_im) : $signed(_GEN_277); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_279 = 5'h1b == _T_12 ? $signed(regsA_15_im) : $signed(_GEN_278); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_281 = 5'h1 == _T_12 ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_282 = 5'h2 == _T_12 ? $signed(regsA_2_re) : $signed(_GEN_281); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_283 = 5'h3 == _T_12 ? $signed(regsA_3_re) : $signed(_GEN_282); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_284 = 5'h4 == _T_12 ? $signed(64'sh0) : $signed(_GEN_283); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_285 = 5'h5 == _T_12 ? $signed(64'sh0) : $signed(_GEN_284); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_286 = 5'h6 == _T_12 ? $signed(64'sh0) : $signed(_GEN_285); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_287 = 5'h7 == _T_12 ? $signed(64'sh0) : $signed(_GEN_286); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_288 = 5'h8 == _T_12 ? $signed(regsA_4_re) : $signed(_GEN_287); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_289 = 5'h9 == _T_12 ? $signed(regsA_5_re) : $signed(_GEN_288); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_290 = 5'ha == _T_12 ? $signed(regsA_6_re) : $signed(_GEN_289); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_291 = 5'hb == _T_12 ? $signed(regsA_7_re) : $signed(_GEN_290); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_292 = 5'hc == _T_12 ? $signed(64'sh0) : $signed(_GEN_291); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_293 = 5'hd == _T_12 ? $signed(64'sh0) : $signed(_GEN_292); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_294 = 5'he == _T_12 ? $signed(64'sh0) : $signed(_GEN_293); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_295 = 5'hf == _T_12 ? $signed(64'sh0) : $signed(_GEN_294); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_296 = 5'h10 == _T_12 ? $signed(regsA_8_re) : $signed(_GEN_295); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_297 = 5'h11 == _T_12 ? $signed(regsA_9_re) : $signed(_GEN_296); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_298 = 5'h12 == _T_12 ? $signed(regsA_10_re) : $signed(_GEN_297); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_299 = 5'h13 == _T_12 ? $signed(regsA_11_re) : $signed(_GEN_298); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_300 = 5'h14 == _T_12 ? $signed(64'sh0) : $signed(_GEN_299); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_301 = 5'h15 == _T_12 ? $signed(64'sh0) : $signed(_GEN_300); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_302 = 5'h16 == _T_12 ? $signed(64'sh0) : $signed(_GEN_301); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_303 = 5'h17 == _T_12 ? $signed(64'sh0) : $signed(_GEN_302); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_304 = 5'h18 == _T_12 ? $signed(regsA_12_re) : $signed(_GEN_303); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_305 = 5'h19 == _T_12 ? $signed(regsA_13_re) : $signed(_GEN_304); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_306 = 5'h1a == _T_12 ? $signed(regsA_14_re) : $signed(_GEN_305); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [63:0] _GEN_307 = 5'h1b == _T_12 ? $signed(regsA_15_re) : $signed(_GEN_306); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [3:0] _T_14 = 1'h0 * 3'h4; // @[Matrix_Mul_V1.scala 162:36]
  wire [4:0] _GEN_329 = {{1'd0}, _T_14}; // @[Matrix_Mul_V1.scala 162:52]
  wire [4:0] _T_16 = _GEN_329 + input_point; // @[Matrix_Mul_V1.scala 162:52]
  wire [63:0] _GEN_317 = 2'h1 == _T_16[1:0] ? $signed(regsB_1_im) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_318 = 2'h2 == _T_16[1:0] ? $signed(regsB_2_im) : $signed(_GEN_317); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_319 = 2'h3 == _T_16[1:0] ? $signed(regsB_3_im) : $signed(_GEN_318); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_321 = 2'h1 == _T_16[1:0] ? $signed(regsB_1_re) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_322 = 2'h2 == _T_16[1:0] ? $signed(regsB_2_re) : $signed(_GEN_321); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [63:0] _GEN_323 = 2'h3 == _T_16[1:0] ? $signed(regsB_3_re) : $signed(_GEN_322); // @[Matrix_Mul_V1.scala 162:{19,19}]
  PE PE ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_clock),
    .io_reset(PE_io_reset),
    .io_in_x_re(PE_io_in_x_re),
    .io_in_x_im(PE_io_in_x_im),
    .io_in_y_re(PE_io_in_y_re),
    .io_in_y_im(PE_io_in_y_im),
    .io_out_pe_re(PE_io_out_pe_re),
    .io_out_pe_im(PE_io_out_pe_im),
    .io_out_x_re(PE_io_out_x_re),
    .io_out_x_im(PE_io_out_x_im),
    .io_out_y_re(PE_io_out_y_re),
    .io_out_y_im(PE_io_out_y_im)
  );
  PE PE_1 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_1_clock),
    .io_reset(PE_1_io_reset),
    .io_in_x_re(PE_1_io_in_x_re),
    .io_in_x_im(PE_1_io_in_x_im),
    .io_in_y_re(PE_1_io_in_y_re),
    .io_in_y_im(PE_1_io_in_y_im),
    .io_out_pe_re(PE_1_io_out_pe_re),
    .io_out_pe_im(PE_1_io_out_pe_im),
    .io_out_x_re(PE_1_io_out_x_re),
    .io_out_x_im(PE_1_io_out_x_im),
    .io_out_y_re(PE_1_io_out_y_re),
    .io_out_y_im(PE_1_io_out_y_im)
  );
  PE PE_2 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_2_clock),
    .io_reset(PE_2_io_reset),
    .io_in_x_re(PE_2_io_in_x_re),
    .io_in_x_im(PE_2_io_in_x_im),
    .io_in_y_re(PE_2_io_in_y_re),
    .io_in_y_im(PE_2_io_in_y_im),
    .io_out_pe_re(PE_2_io_out_pe_re),
    .io_out_pe_im(PE_2_io_out_pe_im),
    .io_out_x_re(PE_2_io_out_x_re),
    .io_out_x_im(PE_2_io_out_x_im),
    .io_out_y_re(PE_2_io_out_y_re),
    .io_out_y_im(PE_2_io_out_y_im)
  );
  PE PE_3 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_3_clock),
    .io_reset(PE_3_io_reset),
    .io_in_x_re(PE_3_io_in_x_re),
    .io_in_x_im(PE_3_io_in_x_im),
    .io_in_y_re(PE_3_io_in_y_re),
    .io_in_y_im(PE_3_io_in_y_im),
    .io_out_pe_re(PE_3_io_out_pe_re),
    .io_out_pe_im(PE_3_io_out_pe_im),
    .io_out_x_re(PE_3_io_out_x_re),
    .io_out_x_im(PE_3_io_out_x_im),
    .io_out_y_re(PE_3_io_out_y_re),
    .io_out_y_im(PE_3_io_out_y_im)
  );
  assign io_matrixC_0_re = PE_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_0_im = PE_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_1_re = PE_1_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_1_im = PE_1_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_2_re = PE_2_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_2_im = PE_2_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_3_re = PE_3_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_3_im = PE_3_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_valid = input_point >= 5'h7; // @[Matrix_Mul_V1.scala 188:20]
  assign PE_clock = clock;
  assign PE_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_io_in_x_re = input_point < 5'h7 ? $signed(_GEN_139) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_io_in_x_im = input_point < 5'h7 ? $signed(_GEN_111) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_io_in_y_re = input_point < 5'h4 ? $signed(_GEN_323) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_io_in_y_im = input_point < 5'h4 ? $signed(_GEN_319) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_1_clock = clock;
  assign PE_1_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_1_io_in_x_re = input_point < 5'h7 ? $signed(_GEN_195) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_1_io_in_x_im = input_point < 5'h7 ? $signed(_GEN_167) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_1_io_in_y_re = PE_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_1_io_in_y_im = PE_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_2_clock = clock;
  assign PE_2_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_2_io_in_x_re = input_point < 5'h7 ? $signed(_GEN_251) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_2_io_in_x_im = input_point < 5'h7 ? $signed(_GEN_223) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_2_io_in_y_re = PE_1_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_2_io_in_y_im = PE_1_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_3_clock = clock;
  assign PE_3_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_3_io_in_x_re = input_point < 5'h7 ? $signed(_GEN_307) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_3_io_in_x_im = input_point < 5'h7 ? $signed(_GEN_279) : $signed(64'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_3_io_in_y_re = PE_2_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_3_io_in_y_im = PE_2_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  always @(posedge clock) begin
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_0_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_0_re <= io_matrixA_0_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_0_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_0_im <= io_matrixA_0_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_1_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_1_re <= io_matrixA_1_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_1_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_1_im <= io_matrixA_1_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_2_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_2_re <= io_matrixA_2_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_2_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_2_im <= io_matrixA_2_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_3_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_3_re <= io_matrixA_3_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_3_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_3_im <= io_matrixA_3_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_4_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_4_re <= io_matrixA_4_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_4_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_4_im <= io_matrixA_4_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_5_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_5_re <= io_matrixA_5_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_5_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_5_im <= io_matrixA_5_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_6_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_6_re <= io_matrixA_6_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_6_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_6_im <= io_matrixA_6_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_7_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_7_re <= io_matrixA_7_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_7_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_7_im <= io_matrixA_7_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_8_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_8_re <= io_matrixA_8_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_8_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_8_im <= io_matrixA_8_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_9_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_9_re <= io_matrixA_9_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_9_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_9_im <= io_matrixA_9_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_10_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_10_re <= io_matrixA_10_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_10_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_10_im <= io_matrixA_10_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_11_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_11_re <= io_matrixA_11_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_11_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_11_im <= io_matrixA_11_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_12_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_12_re <= io_matrixA_12_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_12_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_12_im <= io_matrixA_12_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_13_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_13_re <= io_matrixA_13_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_13_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_13_im <= io_matrixA_13_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_14_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_14_re <= io_matrixA_14_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_14_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_14_im <= io_matrixA_14_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_15_re <= 64'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_15_re <= io_matrixA_15_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_15_im <= 64'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_15_im <= io_matrixA_15_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_0_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_0_re <= io_matrixB_0_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_0_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_0_im <= io_matrixB_0_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_1_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_1_re <= io_matrixB_1_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_1_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_1_im <= io_matrixB_1_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_2_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_2_re <= io_matrixB_2_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_2_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_2_im <= io_matrixB_2_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_3_re <= 64'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_3_re <= io_matrixB_3_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_3_im <= 64'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_3_im <= io_matrixB_3_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      input_point <= 5'h0; // @[Matrix_Mul_V1.scala 99:17]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      input_point <= 5'h0; // @[Matrix_Mul_V1.scala 108:17]
    end else begin
      input_point <= _input_point_T_1; // @[Matrix_Mul_V1.scala 116:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regsA_0_re = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regsA_0_im = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  regsA_1_re = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  regsA_1_im = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  regsA_2_re = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  regsA_2_im = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  regsA_3_re = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  regsA_3_im = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  regsA_4_re = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  regsA_4_im = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  regsA_5_re = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  regsA_5_im = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  regsA_6_re = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  regsA_6_im = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  regsA_7_re = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  regsA_7_im = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  regsA_8_re = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  regsA_8_im = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  regsA_9_re = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  regsA_9_im = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  regsA_10_re = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  regsA_10_im = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  regsA_11_re = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  regsA_11_im = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  regsA_12_re = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  regsA_12_im = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  regsA_13_re = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  regsA_13_im = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  regsA_14_re = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  regsA_14_im = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  regsA_15_re = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  regsA_15_im = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  regsB_0_re = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  regsB_0_im = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  regsB_1_re = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  regsB_1_im = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  regsB_2_re = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  regsB_2_im = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  regsB_3_re = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  regsB_3_im = _RAND_39[63:0];
  _RAND_40 = {1{`RANDOM}};
  input_point = _RAND_40[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module matrix_conjugate(
  input  [63:0] io_matrixIn_0_re,
  input  [63:0] io_matrixIn_0_im,
  input  [63:0] io_matrixIn_1_re,
  input  [63:0] io_matrixIn_1_im,
  input  [63:0] io_matrixIn_2_re,
  input  [63:0] io_matrixIn_2_im,
  input  [63:0] io_matrixIn_3_re,
  input  [63:0] io_matrixIn_3_im,
  output [63:0] io_matrixOut_0_re,
  output [63:0] io_matrixOut_0_im,
  output [63:0] io_matrixOut_1_re,
  output [63:0] io_matrixOut_1_im,
  output [63:0] io_matrixOut_2_re,
  output [63:0] io_matrixOut_2_im,
  output [63:0] io_matrixOut_3_re,
  output [63:0] io_matrixOut_3_im
);
  assign io_matrixOut_0_re = io_matrixIn_0_re; // @[Matrix_Conjugate.scala 22:34]
  assign io_matrixOut_0_im = 64'sh0 - $signed(io_matrixIn_0_im); // @[Matrix_Conjugate.scala 23:37]
  assign io_matrixOut_1_re = io_matrixIn_1_re; // @[Matrix_Conjugate.scala 22:34]
  assign io_matrixOut_1_im = 64'sh0 - $signed(io_matrixIn_1_im); // @[Matrix_Conjugate.scala 23:37]
  assign io_matrixOut_2_re = io_matrixIn_2_re; // @[Matrix_Conjugate.scala 22:34]
  assign io_matrixOut_2_im = 64'sh0 - $signed(io_matrixIn_2_im); // @[Matrix_Conjugate.scala 23:37]
  assign io_matrixOut_3_re = io_matrixIn_3_re; // @[Matrix_Conjugate.scala 22:34]
  assign io_matrixOut_3_im = 64'sh0 - $signed(io_matrixIn_3_im); // @[Matrix_Conjugate.scala 23:37]
endmodule
module matrix_transpose(
  input  [63:0] io_matrixIn_0_re,
  input  [63:0] io_matrixIn_0_im,
  input  [63:0] io_matrixIn_1_re,
  input  [63:0] io_matrixIn_1_im,
  input  [63:0] io_matrixIn_2_re,
  input  [63:0] io_matrixIn_2_im,
  input  [63:0] io_matrixIn_3_re,
  input  [63:0] io_matrixIn_3_im,
  output [63:0] io_matrixOut_0_re,
  output [63:0] io_matrixOut_0_im,
  output [63:0] io_matrixOut_1_re,
  output [63:0] io_matrixOut_1_im,
  output [63:0] io_matrixOut_2_re,
  output [63:0] io_matrixOut_2_im,
  output [63:0] io_matrixOut_3_re,
  output [63:0] io_matrixOut_3_im
);
  assign io_matrixOut_0_re = io_matrixIn_0_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_0_im = io_matrixIn_0_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_1_re = io_matrixIn_1_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_1_im = io_matrixIn_1_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_2_re = io_matrixIn_2_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_2_im = io_matrixIn_2_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_3_re = io_matrixIn_3_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_3_im = io_matrixIn_3_im; // @[Matrix_Transpose.scala 22:31]
endmodule
module matirx_conjugate_transpose(
  input  [63:0] io_matrixIn_0_re,
  input  [63:0] io_matrixIn_0_im,
  input  [63:0] io_matrixIn_1_re,
  input  [63:0] io_matrixIn_1_im,
  input  [63:0] io_matrixIn_2_re,
  input  [63:0] io_matrixIn_2_im,
  input  [63:0] io_matrixIn_3_re,
  input  [63:0] io_matrixIn_3_im,
  output [63:0] io_matrixOut_0_re,
  output [63:0] io_matrixOut_0_im,
  output [63:0] io_matrixOut_1_re,
  output [63:0] io_matrixOut_1_im,
  output [63:0] io_matrixOut_2_re,
  output [63:0] io_matrixOut_2_im,
  output [63:0] io_matrixOut_3_re,
  output [63:0] io_matrixOut_3_im
);
  wire [63:0] unit_io_matrixIn_0_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_0_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_1_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_1_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_2_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_2_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_3_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_3_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_0_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_0_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_1_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_1_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_2_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_2_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_3_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_3_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_1_io_matrixIn_0_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_0_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_1_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_1_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_2_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_2_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_3_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_3_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_0_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_0_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_1_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_1_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_2_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_2_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_3_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_3_im; // @[Matrix_Transpose.scala 36:22]
  matrix_conjugate unit ( // @[Matrix_Conjugate.scala 37:22]
    .io_matrixIn_0_re(unit_io_matrixIn_0_re),
    .io_matrixIn_0_im(unit_io_matrixIn_0_im),
    .io_matrixIn_1_re(unit_io_matrixIn_1_re),
    .io_matrixIn_1_im(unit_io_matrixIn_1_im),
    .io_matrixIn_2_re(unit_io_matrixIn_2_re),
    .io_matrixIn_2_im(unit_io_matrixIn_2_im),
    .io_matrixIn_3_re(unit_io_matrixIn_3_re),
    .io_matrixIn_3_im(unit_io_matrixIn_3_im),
    .io_matrixOut_0_re(unit_io_matrixOut_0_re),
    .io_matrixOut_0_im(unit_io_matrixOut_0_im),
    .io_matrixOut_1_re(unit_io_matrixOut_1_re),
    .io_matrixOut_1_im(unit_io_matrixOut_1_im),
    .io_matrixOut_2_re(unit_io_matrixOut_2_re),
    .io_matrixOut_2_im(unit_io_matrixOut_2_im),
    .io_matrixOut_3_re(unit_io_matrixOut_3_re),
    .io_matrixOut_3_im(unit_io_matrixOut_3_im)
  );
  matrix_transpose unit_1 ( // @[Matrix_Transpose.scala 36:22]
    .io_matrixIn_0_re(unit_1_io_matrixIn_0_re),
    .io_matrixIn_0_im(unit_1_io_matrixIn_0_im),
    .io_matrixIn_1_re(unit_1_io_matrixIn_1_re),
    .io_matrixIn_1_im(unit_1_io_matrixIn_1_im),
    .io_matrixIn_2_re(unit_1_io_matrixIn_2_re),
    .io_matrixIn_2_im(unit_1_io_matrixIn_2_im),
    .io_matrixIn_3_re(unit_1_io_matrixIn_3_re),
    .io_matrixIn_3_im(unit_1_io_matrixIn_3_im),
    .io_matrixOut_0_re(unit_1_io_matrixOut_0_re),
    .io_matrixOut_0_im(unit_1_io_matrixOut_0_im),
    .io_matrixOut_1_re(unit_1_io_matrixOut_1_re),
    .io_matrixOut_1_im(unit_1_io_matrixOut_1_im),
    .io_matrixOut_2_re(unit_1_io_matrixOut_2_re),
    .io_matrixOut_2_im(unit_1_io_matrixOut_2_im),
    .io_matrixOut_3_re(unit_1_io_matrixOut_3_re),
    .io_matrixOut_3_im(unit_1_io_matrixOut_3_im)
  );
  assign io_matrixOut_0_re = unit_1_io_matrixOut_0_re; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_0_im = unit_1_io_matrixOut_0_im; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_1_re = unit_1_io_matrixOut_1_re; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_1_im = unit_1_io_matrixOut_1_im; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_2_re = unit_1_io_matrixOut_2_re; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_2_im = unit_1_io_matrixOut_2_im; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_3_re = unit_1_io_matrixOut_3_re; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_3_im = unit_1_io_matrixOut_3_im; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign unit_io_matrixIn_0_re = io_matrixIn_0_re; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_0_im = io_matrixIn_0_im; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_1_re = io_matrixIn_1_re; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_1_im = io_matrixIn_1_im; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_2_re = io_matrixIn_2_re; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_2_im = io_matrixIn_2_im; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_3_re = io_matrixIn_3_re; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_3_im = io_matrixIn_3_im; // @[Matrix_Conjugate.scala 38:22]
  assign unit_1_io_matrixIn_0_re = unit_io_matrixOut_0_re; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_0_im = unit_io_matrixOut_0_im; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_1_re = unit_io_matrixOut_1_re; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_1_im = unit_io_matrixOut_1_im; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_2_re = unit_io_matrixOut_2_re; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_2_im = unit_io_matrixOut_2_im; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_3_re = unit_io_matrixOut_3_re; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_3_im = unit_io_matrixOut_3_im; // @[Matrix_Transpose.scala 37:22]
endmodule
module optimal_weight_vector(
  input         clock,
  input         reset,
  input         io_reset,
  input         io_ready,
  input  [63:0] io_matrixS_0_re,
  input  [63:0] io_matrixS_0_im,
  input  [63:0] io_matrixS_1_re,
  input  [63:0] io_matrixS_1_im,
  input  [63:0] io_matrixS_2_re,
  input  [63:0] io_matrixS_2_im,
  input  [63:0] io_matrixS_3_re,
  input  [63:0] io_matrixS_3_im,
  input  [63:0] io_matrixR_Inv_0_re,
  input  [63:0] io_matrixR_Inv_0_im,
  input  [63:0] io_matrixR_Inv_1_re,
  input  [63:0] io_matrixR_Inv_1_im,
  input  [63:0] io_matrixR_Inv_2_re,
  input  [63:0] io_matrixR_Inv_2_im,
  input  [63:0] io_matrixR_Inv_3_re,
  input  [63:0] io_matrixR_Inv_3_im,
  input  [63:0] io_matrixR_Inv_4_re,
  input  [63:0] io_matrixR_Inv_4_im,
  input  [63:0] io_matrixR_Inv_5_re,
  input  [63:0] io_matrixR_Inv_5_im,
  input  [63:0] io_matrixR_Inv_6_re,
  input  [63:0] io_matrixR_Inv_6_im,
  input  [63:0] io_matrixR_Inv_7_re,
  input  [63:0] io_matrixR_Inv_7_im,
  input  [63:0] io_matrixR_Inv_8_re,
  input  [63:0] io_matrixR_Inv_8_im,
  input  [63:0] io_matrixR_Inv_9_re,
  input  [63:0] io_matrixR_Inv_9_im,
  input  [63:0] io_matrixR_Inv_10_re,
  input  [63:0] io_matrixR_Inv_10_im,
  input  [63:0] io_matrixR_Inv_11_re,
  input  [63:0] io_matrixR_Inv_11_im,
  input  [63:0] io_matrixR_Inv_12_re,
  input  [63:0] io_matrixR_Inv_12_im,
  input  [63:0] io_matrixR_Inv_13_re,
  input  [63:0] io_matrixR_Inv_13_im,
  input  [63:0] io_matrixR_Inv_14_re,
  input  [63:0] io_matrixR_Inv_14_im,
  input  [63:0] io_matrixR_Inv_15_re,
  input  [63:0] io_matrixR_Inv_15_im,
  output [63:0] io_matrixOut_0_re,
  output [63:0] io_matrixOut_0_im,
  output [63:0] io_matrixOut_1_re,
  output [63:0] io_matrixOut_1_im,
  output [63:0] io_matrixOut_2_re,
  output [63:0] io_matrixOut_2_im,
  output [63:0] io_matrixOut_3_re,
  output [63:0] io_matrixOut_3_im,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [31:0] _RAND_42;
`endif // RANDOMIZE_REG_INIT
  wire  complex_matirx_mul_unit_clock; // @[Optimal_Weight_Vector.scala 38:54]
  wire  complex_matirx_mul_unit_io_reset; // @[Optimal_Weight_Vector.scala 38:54]
  wire  complex_matirx_mul_unit_io_ready; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_0_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_0_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_1_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_1_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_2_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_2_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_3_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_3_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_4_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_4_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_5_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_5_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_6_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_6_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_7_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_7_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_8_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_8_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_9_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_9_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_10_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_10_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_11_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_11_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_12_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_12_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_13_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_13_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_14_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_14_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_15_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixA_15_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixB_0_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixB_0_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixB_1_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixB_1_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixB_2_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixB_2_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixB_3_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixB_3_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_0_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_0_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_1_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_1_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_2_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_2_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_3_re; // @[Optimal_Weight_Vector.scala 38:54]
  wire [63:0] complex_matirx_mul_unit_io_matrixC_3_im; // @[Optimal_Weight_Vector.scala 38:54]
  wire  complex_matirx_mul_unit_io_valid; // @[Optimal_Weight_Vector.scala 38:54]
  wire  complex_divide_unit_clock; // @[Optimal_Weight_Vector.scala 39:58]
  wire  complex_divide_unit_reset; // @[Optimal_Weight_Vector.scala 39:58]
  wire [63:0] complex_divide_unit_io_op2_re; // @[Optimal_Weight_Vector.scala 39:58]
  wire [63:0] complex_divide_unit_io_op2_im; // @[Optimal_Weight_Vector.scala 39:58]
  wire [63:0] complex_divide_unit_io_res_re; // @[Optimal_Weight_Vector.scala 39:58]
  wire [63:0] complex_divide_unit_io_res_im; // @[Optimal_Weight_Vector.scala 39:58]
  wire [63:0] S_c_t_unit_io_matrixIn_0_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] S_c_t_unit_io_matrixIn_0_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] S_c_t_unit_io_matrixIn_1_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] S_c_t_unit_io_matrixIn_1_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] S_c_t_unit_io_matrixIn_2_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] S_c_t_unit_io_matrixIn_2_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] S_c_t_unit_io_matrixIn_3_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] S_c_t_unit_io_matrixIn_3_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] S_c_t_unit_io_matrixOut_0_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] S_c_t_unit_io_matrixOut_0_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] S_c_t_unit_io_matrixOut_1_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] S_c_t_unit_io_matrixOut_1_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] S_c_t_unit_io_matrixOut_2_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] S_c_t_unit_io_matrixOut_2_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] S_c_t_unit_io_matrixOut_3_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] S_c_t_unit_io_matrixOut_3_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] io_matrixOut_0_mul_io_op1_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_0_mul_io_op1_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_0_mul_io_op2_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_0_mul_io_op2_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_0_mul_io_res_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_0_mul_io_res_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_1_mul_io_op1_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_1_mul_io_op1_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_1_mul_io_op2_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_1_mul_io_op2_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_1_mul_io_res_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_1_mul_io_res_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_2_mul_io_op1_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_2_mul_io_op1_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_2_mul_io_op2_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_2_mul_io_op2_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_2_mul_io_res_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_2_mul_io_res_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_3_mul_io_op1_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_3_mul_io_op1_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_3_mul_io_op2_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_3_mul_io_op2_im; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_3_mul_io_res_re; // @[Complex_Operater.scala 47:21]
  wire [63:0] io_matrixOut_3_mul_io_res_im; // @[Complex_Operater.scala 47:21]
  reg [63:0] matrix_R_Comp_0_re; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_0_im; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_1_re; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_1_im; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_2_re; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_2_im; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_3_re; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_3_im; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_4_re; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_4_im; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_5_re; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_5_im; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_6_re; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_6_im; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_7_re; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_7_im; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_8_re; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_8_im; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_9_re; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_9_im; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_10_re; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_10_im; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_11_re; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_11_im; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_12_re; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_12_im; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_13_re; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_13_im; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_14_re; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_14_im; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_15_re; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_R_Comp_15_im; // @[Optimal_Weight_Vector.scala 33:40]
  reg [63:0] matrix_S_Comp_0_re; // @[Optimal_Weight_Vector.scala 34:40]
  reg [63:0] matrix_S_Comp_0_im; // @[Optimal_Weight_Vector.scala 34:40]
  reg [63:0] matrix_S_Comp_1_re; // @[Optimal_Weight_Vector.scala 34:40]
  reg [63:0] matrix_S_Comp_1_im; // @[Optimal_Weight_Vector.scala 34:40]
  reg [63:0] matrix_S_Comp_2_re; // @[Optimal_Weight_Vector.scala 34:40]
  reg [63:0] matrix_S_Comp_2_im; // @[Optimal_Weight_Vector.scala 34:40]
  reg [63:0] matrix_S_Comp_3_re; // @[Optimal_Weight_Vector.scala 34:40]
  reg [63:0] matrix_S_Comp_3_im; // @[Optimal_Weight_Vector.scala 34:40]
  reg [63:0] u_re; // @[Optimal_Weight_Vector.scala 35:23]
  reg [63:0] u_im; // @[Optimal_Weight_Vector.scala 35:23]
  reg [7:0] status; // @[Optimal_Weight_Vector.scala 36:29]
  wire [7:0] _status_T_1 = status + 8'h1; // @[Optimal_Weight_Vector.scala 80:24]
  wire [63:0] _GEN_0 = complex_matirx_mul_unit_io_valid ? $signed(complex_matirx_mul_unit_io_matrixC_0_im) : $signed(
    matrix_R_Comp_0_im); // @[Optimal_Weight_Vector.scala 84:46 86:28 33:40]
  wire [63:0] _GEN_1 = complex_matirx_mul_unit_io_valid ? $signed(complex_matirx_mul_unit_io_matrixC_0_re) : $signed(
    matrix_R_Comp_0_re); // @[Optimal_Weight_Vector.scala 84:46 86:28 33:40]
  wire [63:0] _GEN_2 = complex_matirx_mul_unit_io_valid ? $signed(complex_matirx_mul_unit_io_matrixC_1_im) : $signed(
    matrix_R_Comp_1_im); // @[Optimal_Weight_Vector.scala 84:46 86:28 33:40]
  wire [63:0] _GEN_3 = complex_matirx_mul_unit_io_valid ? $signed(complex_matirx_mul_unit_io_matrixC_1_re) : $signed(
    matrix_R_Comp_1_re); // @[Optimal_Weight_Vector.scala 84:46 86:28 33:40]
  wire [63:0] _GEN_4 = complex_matirx_mul_unit_io_valid ? $signed(complex_matirx_mul_unit_io_matrixC_2_im) : $signed(
    matrix_R_Comp_2_im); // @[Optimal_Weight_Vector.scala 84:46 86:28 33:40]
  wire [63:0] _GEN_5 = complex_matirx_mul_unit_io_valid ? $signed(complex_matirx_mul_unit_io_matrixC_2_re) : $signed(
    matrix_R_Comp_2_re); // @[Optimal_Weight_Vector.scala 84:46 86:28 33:40]
  wire [63:0] _GEN_6 = complex_matirx_mul_unit_io_valid ? $signed(complex_matirx_mul_unit_io_matrixC_3_im) : $signed(
    matrix_R_Comp_3_im); // @[Optimal_Weight_Vector.scala 84:46 86:28 33:40]
  wire [63:0] _GEN_7 = complex_matirx_mul_unit_io_valid ? $signed(complex_matirx_mul_unit_io_matrixC_3_re) : $signed(
    matrix_R_Comp_3_re); // @[Optimal_Weight_Vector.scala 84:46 86:28 33:40]
  wire [7:0] _GEN_8 = complex_matirx_mul_unit_io_valid ? _status_T_1 : status; // @[Optimal_Weight_Vector.scala 84:46 88:16 36:29]
  wire  _T_2 = status == 8'h3; // @[Optimal_Weight_Vector.scala 90:23]
  wire [63:0] _GEN_9 = complex_matirx_mul_unit_io_valid ? $signed(complex_matirx_mul_unit_io_matrixC_0_im) : $signed(
    u_im); // @[Optimal_Weight_Vector.scala 103:46 104:11 35:23]
  wire [63:0] _GEN_10 = complex_matirx_mul_unit_io_valid ? $signed(complex_matirx_mul_unit_io_matrixC_0_re) : $signed(
    u_re); // @[Optimal_Weight_Vector.scala 103:46 104:11 35:23]
  wire [63:0] _GEN_12 = status <= 8'h32 ? $signed(u_im) : $signed(64'sh100000000); // @[Optimal_Weight_Vector.scala 107:54 109:34 47:33]
  wire [63:0] _GEN_13 = status <= 8'h32 ? $signed(u_re) : $signed(64'sh100000000); // @[Optimal_Weight_Vector.scala 107:54 109:34 46:33]
  wire [7:0] _GEN_14 = status <= 8'h32 ? _status_T_1 : status; // @[Optimal_Weight_Vector.scala 107:54 110:14 36:29]
  wire [63:0] _GEN_16 = status == 8'h4 ? $signed(_GEN_9) : $signed(u_im); // @[Optimal_Weight_Vector.scala 100:32 35:23]
  wire [63:0] _GEN_17 = status == 8'h4 ? $signed(_GEN_10) : $signed(u_re); // @[Optimal_Weight_Vector.scala 100:32 35:23]
  wire [7:0] _GEN_18 = status == 8'h4 ? _GEN_8 : _GEN_14; // @[Optimal_Weight_Vector.scala 100:32]
  wire [63:0] _GEN_19 = status == 8'h4 ? $signed(64'sh100000000) : $signed(_GEN_12); // @[Optimal_Weight_Vector.scala 100:32 47:33]
  wire [63:0] _GEN_20 = status == 8'h4 ? $signed(64'sh100000000) : $signed(_GEN_13); // @[Optimal_Weight_Vector.scala 100:32 46:33]
  wire [63:0] _GEN_22 = S_c_t_unit_io_matrixOut_0_im; // @[Optimal_Weight_Vector.scala 90:32 96:47]
  wire [63:0] _GEN_23 = S_c_t_unit_io_matrixOut_0_re; // @[Optimal_Weight_Vector.scala 90:32 96:47]
  wire [63:0] _GEN_26 = S_c_t_unit_io_matrixOut_1_im; // @[Optimal_Weight_Vector.scala 90:32 96:47]
  wire [63:0] _GEN_27 = S_c_t_unit_io_matrixOut_1_re; // @[Optimal_Weight_Vector.scala 90:32 96:47]
  wire [63:0] _GEN_30 = S_c_t_unit_io_matrixOut_2_im; // @[Optimal_Weight_Vector.scala 90:32 96:47]
  wire [63:0] _GEN_31 = S_c_t_unit_io_matrixOut_2_re; // @[Optimal_Weight_Vector.scala 90:32 96:47]
  wire [63:0] _GEN_34 = S_c_t_unit_io_matrixOut_3_im; // @[Optimal_Weight_Vector.scala 90:32 96:47]
  wire [63:0] _GEN_35 = S_c_t_unit_io_matrixOut_3_re; // @[Optimal_Weight_Vector.scala 90:32 96:47]
  wire [7:0] _GEN_38 = status == 8'h3 ? _status_T_1 : _GEN_18; // @[Optimal_Weight_Vector.scala 90:32 99:14]
  wire [63:0] _GEN_39 = status == 8'h3 ? $signed(u_im) : $signed(_GEN_16); // @[Optimal_Weight_Vector.scala 35:23 90:32]
  wire [63:0] _GEN_40 = status == 8'h3 ? $signed(u_re) : $signed(_GEN_17); // @[Optimal_Weight_Vector.scala 35:23 90:32]
  wire [63:0] _GEN_41 = status == 8'h3 ? $signed(64'sh100000000) : $signed(_GEN_19); // @[Optimal_Weight_Vector.scala 90:32 47:33]
  wire [63:0] _GEN_42 = status == 8'h3 ? $signed(64'sh100000000) : $signed(_GEN_20); // @[Optimal_Weight_Vector.scala 90:32 46:33]
  wire  _GEN_43 = status == 8'h2 ? 1'h0 : _T_2; // @[Optimal_Weight_Vector.scala 81:32 83:40]
  wire [7:0] _GEN_52 = status == 8'h2 ? _GEN_8 : _GEN_38; // @[Optimal_Weight_Vector.scala 81:32]
  wire [63:0] _GEN_71 = status == 8'h2 ? $signed(64'sh100000000) : $signed(_GEN_41); // @[Optimal_Weight_Vector.scala 81:32 47:33]
  wire [63:0] _GEN_72 = status == 8'h2 ? $signed(64'sh100000000) : $signed(_GEN_42); // @[Optimal_Weight_Vector.scala 81:32 46:33]
  wire [63:0] _GEN_125 = status == 8'h1 ? $signed(64'sh100000000) : $signed(_GEN_71); // @[Optimal_Weight_Vector.scala 75:26 47:33]
  wire [63:0] _GEN_126 = status == 8'h1 ? $signed(64'sh100000000) : $signed(_GEN_72); // @[Optimal_Weight_Vector.scala 75:26 46:33]
  wire [63:0] _GEN_211 = io_ready ? $signed(64'sh100000000) : $signed(_GEN_125); // @[Optimal_Weight_Vector.scala 69:24 47:33]
  wire [63:0] _GEN_212 = io_ready ? $signed(64'sh100000000) : $signed(_GEN_126); // @[Optimal_Weight_Vector.scala 69:24 46:33]
  matrix_mul_v1_3 complex_matirx_mul_unit ( // @[Optimal_Weight_Vector.scala 38:54]
    .clock(complex_matirx_mul_unit_clock),
    .io_reset(complex_matirx_mul_unit_io_reset),
    .io_ready(complex_matirx_mul_unit_io_ready),
    .io_matrixA_0_re(complex_matirx_mul_unit_io_matrixA_0_re),
    .io_matrixA_0_im(complex_matirx_mul_unit_io_matrixA_0_im),
    .io_matrixA_1_re(complex_matirx_mul_unit_io_matrixA_1_re),
    .io_matrixA_1_im(complex_matirx_mul_unit_io_matrixA_1_im),
    .io_matrixA_2_re(complex_matirx_mul_unit_io_matrixA_2_re),
    .io_matrixA_2_im(complex_matirx_mul_unit_io_matrixA_2_im),
    .io_matrixA_3_re(complex_matirx_mul_unit_io_matrixA_3_re),
    .io_matrixA_3_im(complex_matirx_mul_unit_io_matrixA_3_im),
    .io_matrixA_4_re(complex_matirx_mul_unit_io_matrixA_4_re),
    .io_matrixA_4_im(complex_matirx_mul_unit_io_matrixA_4_im),
    .io_matrixA_5_re(complex_matirx_mul_unit_io_matrixA_5_re),
    .io_matrixA_5_im(complex_matirx_mul_unit_io_matrixA_5_im),
    .io_matrixA_6_re(complex_matirx_mul_unit_io_matrixA_6_re),
    .io_matrixA_6_im(complex_matirx_mul_unit_io_matrixA_6_im),
    .io_matrixA_7_re(complex_matirx_mul_unit_io_matrixA_7_re),
    .io_matrixA_7_im(complex_matirx_mul_unit_io_matrixA_7_im),
    .io_matrixA_8_re(complex_matirx_mul_unit_io_matrixA_8_re),
    .io_matrixA_8_im(complex_matirx_mul_unit_io_matrixA_8_im),
    .io_matrixA_9_re(complex_matirx_mul_unit_io_matrixA_9_re),
    .io_matrixA_9_im(complex_matirx_mul_unit_io_matrixA_9_im),
    .io_matrixA_10_re(complex_matirx_mul_unit_io_matrixA_10_re),
    .io_matrixA_10_im(complex_matirx_mul_unit_io_matrixA_10_im),
    .io_matrixA_11_re(complex_matirx_mul_unit_io_matrixA_11_re),
    .io_matrixA_11_im(complex_matirx_mul_unit_io_matrixA_11_im),
    .io_matrixA_12_re(complex_matirx_mul_unit_io_matrixA_12_re),
    .io_matrixA_12_im(complex_matirx_mul_unit_io_matrixA_12_im),
    .io_matrixA_13_re(complex_matirx_mul_unit_io_matrixA_13_re),
    .io_matrixA_13_im(complex_matirx_mul_unit_io_matrixA_13_im),
    .io_matrixA_14_re(complex_matirx_mul_unit_io_matrixA_14_re),
    .io_matrixA_14_im(complex_matirx_mul_unit_io_matrixA_14_im),
    .io_matrixA_15_re(complex_matirx_mul_unit_io_matrixA_15_re),
    .io_matrixA_15_im(complex_matirx_mul_unit_io_matrixA_15_im),
    .io_matrixB_0_re(complex_matirx_mul_unit_io_matrixB_0_re),
    .io_matrixB_0_im(complex_matirx_mul_unit_io_matrixB_0_im),
    .io_matrixB_1_re(complex_matirx_mul_unit_io_matrixB_1_re),
    .io_matrixB_1_im(complex_matirx_mul_unit_io_matrixB_1_im),
    .io_matrixB_2_re(complex_matirx_mul_unit_io_matrixB_2_re),
    .io_matrixB_2_im(complex_matirx_mul_unit_io_matrixB_2_im),
    .io_matrixB_3_re(complex_matirx_mul_unit_io_matrixB_3_re),
    .io_matrixB_3_im(complex_matirx_mul_unit_io_matrixB_3_im),
    .io_matrixC_0_re(complex_matirx_mul_unit_io_matrixC_0_re),
    .io_matrixC_0_im(complex_matirx_mul_unit_io_matrixC_0_im),
    .io_matrixC_1_re(complex_matirx_mul_unit_io_matrixC_1_re),
    .io_matrixC_1_im(complex_matirx_mul_unit_io_matrixC_1_im),
    .io_matrixC_2_re(complex_matirx_mul_unit_io_matrixC_2_re),
    .io_matrixC_2_im(complex_matirx_mul_unit_io_matrixC_2_im),
    .io_matrixC_3_re(complex_matirx_mul_unit_io_matrixC_3_re),
    .io_matrixC_3_im(complex_matirx_mul_unit_io_matrixC_3_im),
    .io_valid(complex_matirx_mul_unit_io_valid)
  );
  cordic_complex_divide complex_divide_unit ( // @[Optimal_Weight_Vector.scala 39:58]
    .clock(complex_divide_unit_clock),
    .reset(complex_divide_unit_reset),
    .io_op2_re(complex_divide_unit_io_op2_re),
    .io_op2_im(complex_divide_unit_io_op2_im),
    .io_res_re(complex_divide_unit_io_res_re),
    .io_res_im(complex_divide_unit_io_res_im)
  );
  matirx_conjugate_transpose S_c_t_unit ( // @[Matirx_Conjugate_Transpose.scala 32:22]
    .io_matrixIn_0_re(S_c_t_unit_io_matrixIn_0_re),
    .io_matrixIn_0_im(S_c_t_unit_io_matrixIn_0_im),
    .io_matrixIn_1_re(S_c_t_unit_io_matrixIn_1_re),
    .io_matrixIn_1_im(S_c_t_unit_io_matrixIn_1_im),
    .io_matrixIn_2_re(S_c_t_unit_io_matrixIn_2_re),
    .io_matrixIn_2_im(S_c_t_unit_io_matrixIn_2_im),
    .io_matrixIn_3_re(S_c_t_unit_io_matrixIn_3_re),
    .io_matrixIn_3_im(S_c_t_unit_io_matrixIn_3_im),
    .io_matrixOut_0_re(S_c_t_unit_io_matrixOut_0_re),
    .io_matrixOut_0_im(S_c_t_unit_io_matrixOut_0_im),
    .io_matrixOut_1_re(S_c_t_unit_io_matrixOut_1_re),
    .io_matrixOut_1_im(S_c_t_unit_io_matrixOut_1_im),
    .io_matrixOut_2_re(S_c_t_unit_io_matrixOut_2_re),
    .io_matrixOut_2_im(S_c_t_unit_io_matrixOut_2_im),
    .io_matrixOut_3_re(S_c_t_unit_io_matrixOut_3_re),
    .io_matrixOut_3_im(S_c_t_unit_io_matrixOut_3_im)
  );
  ComplexMul io_matrixOut_0_mul ( // @[Complex_Operater.scala 47:21]
    .io_op1_re(io_matrixOut_0_mul_io_op1_re),
    .io_op1_im(io_matrixOut_0_mul_io_op1_im),
    .io_op2_re(io_matrixOut_0_mul_io_op2_re),
    .io_op2_im(io_matrixOut_0_mul_io_op2_im),
    .io_res_re(io_matrixOut_0_mul_io_res_re),
    .io_res_im(io_matrixOut_0_mul_io_res_im)
  );
  ComplexMul io_matrixOut_1_mul ( // @[Complex_Operater.scala 47:21]
    .io_op1_re(io_matrixOut_1_mul_io_op1_re),
    .io_op1_im(io_matrixOut_1_mul_io_op1_im),
    .io_op2_re(io_matrixOut_1_mul_io_op2_re),
    .io_op2_im(io_matrixOut_1_mul_io_op2_im),
    .io_res_re(io_matrixOut_1_mul_io_res_re),
    .io_res_im(io_matrixOut_1_mul_io_res_im)
  );
  ComplexMul io_matrixOut_2_mul ( // @[Complex_Operater.scala 47:21]
    .io_op1_re(io_matrixOut_2_mul_io_op1_re),
    .io_op1_im(io_matrixOut_2_mul_io_op1_im),
    .io_op2_re(io_matrixOut_2_mul_io_op2_re),
    .io_op2_im(io_matrixOut_2_mul_io_op2_im),
    .io_res_re(io_matrixOut_2_mul_io_res_re),
    .io_res_im(io_matrixOut_2_mul_io_res_im)
  );
  ComplexMul io_matrixOut_3_mul ( // @[Complex_Operater.scala 47:21]
    .io_op1_re(io_matrixOut_3_mul_io_op1_re),
    .io_op1_im(io_matrixOut_3_mul_io_op1_im),
    .io_op2_re(io_matrixOut_3_mul_io_op2_re),
    .io_op2_im(io_matrixOut_3_mul_io_op2_im),
    .io_res_re(io_matrixOut_3_mul_io_res_re),
    .io_res_im(io_matrixOut_3_mul_io_res_im)
  );
  assign io_matrixOut_0_re = io_matrixOut_0_mul_io_res_re; // @[Optimal_Weight_Vector.scala 121:21]
  assign io_matrixOut_0_im = io_matrixOut_0_mul_io_res_im; // @[Optimal_Weight_Vector.scala 121:21]
  assign io_matrixOut_1_re = io_matrixOut_1_mul_io_res_re; // @[Optimal_Weight_Vector.scala 121:21]
  assign io_matrixOut_1_im = io_matrixOut_1_mul_io_res_im; // @[Optimal_Weight_Vector.scala 121:21]
  assign io_matrixOut_2_re = io_matrixOut_2_mul_io_res_re; // @[Optimal_Weight_Vector.scala 121:21]
  assign io_matrixOut_2_im = io_matrixOut_2_mul_io_res_im; // @[Optimal_Weight_Vector.scala 121:21]
  assign io_matrixOut_3_re = io_matrixOut_3_mul_io_res_re; // @[Optimal_Weight_Vector.scala 121:21]
  assign io_matrixOut_3_im = io_matrixOut_3_mul_io_res_im; // @[Optimal_Weight_Vector.scala 121:21]
  assign io_valid = status > 8'h32; // @[Optimal_Weight_Vector.scala 114:15]
  assign complex_matirx_mul_unit_clock = clock;
  assign complex_matirx_mul_unit_io_reset = io_reset; // @[Optimal_Weight_Vector.scala 40:36]
  assign complex_matirx_mul_unit_io_ready = status == 8'h1 | _GEN_43; // @[Optimal_Weight_Vector.scala 75:26 77:40]
  assign complex_matirx_mul_unit_io_matrixA_0_re = status == 8'h1 ? $signed(matrix_R_Comp_0_re) : $signed(_GEN_23); // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_0_im = status == 8'h1 ? $signed(matrix_R_Comp_0_im) : $signed(_GEN_22); // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_1_re = status == 8'h1 ? $signed(matrix_R_Comp_1_re) : $signed(_GEN_27); // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_1_im = status == 8'h1 ? $signed(matrix_R_Comp_1_im) : $signed(_GEN_26); // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_2_re = status == 8'h1 ? $signed(matrix_R_Comp_2_re) : $signed(_GEN_31); // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_2_im = status == 8'h1 ? $signed(matrix_R_Comp_2_im) : $signed(_GEN_30); // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_3_re = status == 8'h1 ? $signed(matrix_R_Comp_3_re) : $signed(_GEN_35); // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_3_im = status == 8'h1 ? $signed(matrix_R_Comp_3_im) : $signed(_GEN_34); // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_4_re = matrix_R_Comp_4_re; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_4_im = matrix_R_Comp_4_im; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_5_re = matrix_R_Comp_5_re; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_5_im = matrix_R_Comp_5_im; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_6_re = matrix_R_Comp_6_re; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_6_im = matrix_R_Comp_6_im; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_7_re = matrix_R_Comp_7_re; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_7_im = matrix_R_Comp_7_im; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_8_re = matrix_R_Comp_8_re; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_8_im = matrix_R_Comp_8_im; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_9_re = matrix_R_Comp_9_re; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_9_im = matrix_R_Comp_9_im; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_10_re = matrix_R_Comp_10_re; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_10_im = matrix_R_Comp_10_im; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_11_re = matrix_R_Comp_11_re; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_11_im = matrix_R_Comp_11_im; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_12_re = matrix_R_Comp_12_re; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_12_im = matrix_R_Comp_12_im; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_13_re = matrix_R_Comp_13_re; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_13_im = matrix_R_Comp_13_im; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_14_re = matrix_R_Comp_14_re; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_14_im = matrix_R_Comp_14_im; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_15_re = matrix_R_Comp_15_re; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixA_15_im = matrix_R_Comp_15_im; // @[Optimal_Weight_Vector.scala 75:26 78:42]
  assign complex_matirx_mul_unit_io_matrixB_0_re = status == 8'h1 ? $signed(matrix_S_Comp_0_re) : $signed(
    matrix_R_Comp_0_re); // @[Optimal_Weight_Vector.scala 75:26 79:42]
  assign complex_matirx_mul_unit_io_matrixB_0_im = status == 8'h1 ? $signed(matrix_S_Comp_0_im) : $signed(
    matrix_R_Comp_0_im); // @[Optimal_Weight_Vector.scala 75:26 79:42]
  assign complex_matirx_mul_unit_io_matrixB_1_re = status == 8'h1 ? $signed(matrix_S_Comp_1_re) : $signed(
    matrix_R_Comp_1_re); // @[Optimal_Weight_Vector.scala 75:26 79:42]
  assign complex_matirx_mul_unit_io_matrixB_1_im = status == 8'h1 ? $signed(matrix_S_Comp_1_im) : $signed(
    matrix_R_Comp_1_im); // @[Optimal_Weight_Vector.scala 75:26 79:42]
  assign complex_matirx_mul_unit_io_matrixB_2_re = status == 8'h1 ? $signed(matrix_S_Comp_2_re) : $signed(
    matrix_R_Comp_2_re); // @[Optimal_Weight_Vector.scala 75:26 79:42]
  assign complex_matirx_mul_unit_io_matrixB_2_im = status == 8'h1 ? $signed(matrix_S_Comp_2_im) : $signed(
    matrix_R_Comp_2_im); // @[Optimal_Weight_Vector.scala 75:26 79:42]
  assign complex_matirx_mul_unit_io_matrixB_3_re = status == 8'h1 ? $signed(matrix_S_Comp_3_re) : $signed(
    matrix_R_Comp_3_re); // @[Optimal_Weight_Vector.scala 75:26 79:42]
  assign complex_matirx_mul_unit_io_matrixB_3_im = status == 8'h1 ? $signed(matrix_S_Comp_3_im) : $signed(
    matrix_R_Comp_3_im); // @[Optimal_Weight_Vector.scala 75:26 79:42]
  assign complex_divide_unit_clock = clock;
  assign complex_divide_unit_reset = reset;
  assign complex_divide_unit_io_op2_re = io_reset ? $signed(64'sh100000000) : $signed(_GEN_212); // @[Optimal_Weight_Vector.scala 56:18 46:33]
  assign complex_divide_unit_io_op2_im = io_reset ? $signed(64'sh100000000) : $signed(_GEN_211); // @[Optimal_Weight_Vector.scala 56:18 47:33]
  assign S_c_t_unit_io_matrixIn_0_re = matrix_S_Comp_0_re; // @[Matirx_Conjugate_Transpose.scala 33:22]
  assign S_c_t_unit_io_matrixIn_0_im = matrix_S_Comp_0_im; // @[Matirx_Conjugate_Transpose.scala 33:22]
  assign S_c_t_unit_io_matrixIn_1_re = matrix_S_Comp_1_re; // @[Matirx_Conjugate_Transpose.scala 33:22]
  assign S_c_t_unit_io_matrixIn_1_im = matrix_S_Comp_1_im; // @[Matirx_Conjugate_Transpose.scala 33:22]
  assign S_c_t_unit_io_matrixIn_2_re = matrix_S_Comp_2_re; // @[Matirx_Conjugate_Transpose.scala 33:22]
  assign S_c_t_unit_io_matrixIn_2_im = matrix_S_Comp_2_im; // @[Matirx_Conjugate_Transpose.scala 33:22]
  assign S_c_t_unit_io_matrixIn_3_re = matrix_S_Comp_3_re; // @[Matirx_Conjugate_Transpose.scala 33:22]
  assign S_c_t_unit_io_matrixIn_3_im = matrix_S_Comp_3_im; // @[Matirx_Conjugate_Transpose.scala 33:22]
  assign io_matrixOut_0_mul_io_op1_re = complex_divide_unit_io_res_re; // @[Complex_Operater.scala 48:16]
  assign io_matrixOut_0_mul_io_op1_im = complex_divide_unit_io_res_im; // @[Complex_Operater.scala 48:16]
  assign io_matrixOut_0_mul_io_op2_re = matrix_R_Comp_0_re; // @[Complex_Operater.scala 49:16]
  assign io_matrixOut_0_mul_io_op2_im = matrix_R_Comp_0_im; // @[Complex_Operater.scala 49:16]
  assign io_matrixOut_1_mul_io_op1_re = complex_divide_unit_io_res_re; // @[Complex_Operater.scala 48:16]
  assign io_matrixOut_1_mul_io_op1_im = complex_divide_unit_io_res_im; // @[Complex_Operater.scala 48:16]
  assign io_matrixOut_1_mul_io_op2_re = matrix_R_Comp_1_re; // @[Complex_Operater.scala 49:16]
  assign io_matrixOut_1_mul_io_op2_im = matrix_R_Comp_1_im; // @[Complex_Operater.scala 49:16]
  assign io_matrixOut_2_mul_io_op1_re = complex_divide_unit_io_res_re; // @[Complex_Operater.scala 48:16]
  assign io_matrixOut_2_mul_io_op1_im = complex_divide_unit_io_res_im; // @[Complex_Operater.scala 48:16]
  assign io_matrixOut_2_mul_io_op2_re = matrix_R_Comp_2_re; // @[Complex_Operater.scala 49:16]
  assign io_matrixOut_2_mul_io_op2_im = matrix_R_Comp_2_im; // @[Complex_Operater.scala 49:16]
  assign io_matrixOut_3_mul_io_op1_re = complex_divide_unit_io_res_re; // @[Complex_Operater.scala 48:16]
  assign io_matrixOut_3_mul_io_op1_im = complex_divide_unit_io_res_im; // @[Complex_Operater.scala 48:16]
  assign io_matrixOut_3_mul_io_op2_re = matrix_R_Comp_3_re; // @[Complex_Operater.scala 49:16]
  assign io_matrixOut_3_mul_io_op2_im = matrix_R_Comp_3_im; // @[Complex_Operater.scala 49:16]
  always @(posedge clock) begin
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_0_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 59:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_0_re <= io_matrixR_Inv_0_re; // @[Optimal_Weight_Vector.scala 71:19]
    end else if (!(status == 8'h1)) begin // @[Optimal_Weight_Vector.scala 75:26]
      if (status == 8'h2) begin // @[Optimal_Weight_Vector.scala 81:32]
        matrix_R_Comp_0_re <= _GEN_1;
      end
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_0_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 60:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_0_im <= io_matrixR_Inv_0_im; // @[Optimal_Weight_Vector.scala 71:19]
    end else if (!(status == 8'h1)) begin // @[Optimal_Weight_Vector.scala 75:26]
      if (status == 8'h2) begin // @[Optimal_Weight_Vector.scala 81:32]
        matrix_R_Comp_0_im <= _GEN_0;
      end
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_1_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 59:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_1_re <= io_matrixR_Inv_1_re; // @[Optimal_Weight_Vector.scala 71:19]
    end else if (!(status == 8'h1)) begin // @[Optimal_Weight_Vector.scala 75:26]
      if (status == 8'h2) begin // @[Optimal_Weight_Vector.scala 81:32]
        matrix_R_Comp_1_re <= _GEN_3;
      end
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_1_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 60:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_1_im <= io_matrixR_Inv_1_im; // @[Optimal_Weight_Vector.scala 71:19]
    end else if (!(status == 8'h1)) begin // @[Optimal_Weight_Vector.scala 75:26]
      if (status == 8'h2) begin // @[Optimal_Weight_Vector.scala 81:32]
        matrix_R_Comp_1_im <= _GEN_2;
      end
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_2_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 59:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_2_re <= io_matrixR_Inv_2_re; // @[Optimal_Weight_Vector.scala 71:19]
    end else if (!(status == 8'h1)) begin // @[Optimal_Weight_Vector.scala 75:26]
      if (status == 8'h2) begin // @[Optimal_Weight_Vector.scala 81:32]
        matrix_R_Comp_2_re <= _GEN_5;
      end
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_2_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 60:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_2_im <= io_matrixR_Inv_2_im; // @[Optimal_Weight_Vector.scala 71:19]
    end else if (!(status == 8'h1)) begin // @[Optimal_Weight_Vector.scala 75:26]
      if (status == 8'h2) begin // @[Optimal_Weight_Vector.scala 81:32]
        matrix_R_Comp_2_im <= _GEN_4;
      end
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_3_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 59:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_3_re <= io_matrixR_Inv_3_re; // @[Optimal_Weight_Vector.scala 71:19]
    end else if (!(status == 8'h1)) begin // @[Optimal_Weight_Vector.scala 75:26]
      if (status == 8'h2) begin // @[Optimal_Weight_Vector.scala 81:32]
        matrix_R_Comp_3_re <= _GEN_7;
      end
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_3_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 60:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_3_im <= io_matrixR_Inv_3_im; // @[Optimal_Weight_Vector.scala 71:19]
    end else if (!(status == 8'h1)) begin // @[Optimal_Weight_Vector.scala 75:26]
      if (status == 8'h2) begin // @[Optimal_Weight_Vector.scala 81:32]
        matrix_R_Comp_3_im <= _GEN_6;
      end
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_4_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 59:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_4_re <= io_matrixR_Inv_4_re; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_4_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 60:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_4_im <= io_matrixR_Inv_4_im; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_5_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 59:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_5_re <= io_matrixR_Inv_5_re; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_5_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 60:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_5_im <= io_matrixR_Inv_5_im; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_6_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 59:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_6_re <= io_matrixR_Inv_6_re; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_6_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 60:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_6_im <= io_matrixR_Inv_6_im; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_7_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 59:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_7_re <= io_matrixR_Inv_7_re; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_7_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 60:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_7_im <= io_matrixR_Inv_7_im; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_8_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 59:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_8_re <= io_matrixR_Inv_8_re; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_8_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 60:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_8_im <= io_matrixR_Inv_8_im; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_9_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 59:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_9_re <= io_matrixR_Inv_9_re; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_9_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 60:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_9_im <= io_matrixR_Inv_9_im; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_10_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 59:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_10_re <= io_matrixR_Inv_10_re; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_10_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 60:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_10_im <= io_matrixR_Inv_10_im; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_11_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 59:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_11_re <= io_matrixR_Inv_11_re; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_11_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 60:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_11_im <= io_matrixR_Inv_11_im; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_12_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 59:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_12_re <= io_matrixR_Inv_12_re; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_12_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 60:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_12_im <= io_matrixR_Inv_12_im; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_13_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 59:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_13_re <= io_matrixR_Inv_13_re; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_13_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 60:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_13_im <= io_matrixR_Inv_13_im; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_14_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 59:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_14_re <= io_matrixR_Inv_14_re; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_14_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 60:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_14_im <= io_matrixR_Inv_14_im; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_15_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 59:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_15_re <= io_matrixR_Inv_15_re; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_R_Comp_15_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 60:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_R_Comp_15_im <= io_matrixR_Inv_15_im; // @[Optimal_Weight_Vector.scala 71:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_S_Comp_0_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 63:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_S_Comp_0_re <= io_matrixS_0_re; // @[Optimal_Weight_Vector.scala 72:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_S_Comp_0_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 64:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_S_Comp_0_im <= io_matrixS_0_im; // @[Optimal_Weight_Vector.scala 72:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_S_Comp_1_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 63:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_S_Comp_1_re <= io_matrixS_1_re; // @[Optimal_Weight_Vector.scala 72:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_S_Comp_1_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 64:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_S_Comp_1_im <= io_matrixS_1_im; // @[Optimal_Weight_Vector.scala 72:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_S_Comp_2_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 63:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_S_Comp_2_re <= io_matrixS_2_re; // @[Optimal_Weight_Vector.scala 72:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_S_Comp_2_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 64:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_S_Comp_2_im <= io_matrixS_2_im; // @[Optimal_Weight_Vector.scala 72:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_S_Comp_3_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 63:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_S_Comp_3_re <= io_matrixS_3_re; // @[Optimal_Weight_Vector.scala 72:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      matrix_S_Comp_3_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 64:27]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      matrix_S_Comp_3_im <= io_matrixS_3_im; // @[Optimal_Weight_Vector.scala 72:19]
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      u_re <= 64'sh0; // @[Optimal_Weight_Vector.scala 66:10]
    end else if (!(io_ready)) begin // @[Optimal_Weight_Vector.scala 69:24]
      if (!(status == 8'h1)) begin // @[Optimal_Weight_Vector.scala 75:26]
        if (!(status == 8'h2)) begin // @[Optimal_Weight_Vector.scala 81:32]
          u_re <= _GEN_40;
        end
      end
    end
    if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      u_im <= 64'sh0; // @[Optimal_Weight_Vector.scala 67:10]
    end else if (!(io_ready)) begin // @[Optimal_Weight_Vector.scala 69:24]
      if (!(status == 8'h1)) begin // @[Optimal_Weight_Vector.scala 75:26]
        if (!(status == 8'h2)) begin // @[Optimal_Weight_Vector.scala 81:32]
          u_im <= _GEN_39;
        end
      end
    end
    if (reset) begin // @[Optimal_Weight_Vector.scala 36:29]
      status <= 8'h0; // @[Optimal_Weight_Vector.scala 36:29]
    end else if (io_reset) begin // @[Optimal_Weight_Vector.scala 56:18]
      status <= 8'h0; // @[Optimal_Weight_Vector.scala 68:12]
    end else if (io_ready) begin // @[Optimal_Weight_Vector.scala 69:24]
      status <= 8'h1; // @[Optimal_Weight_Vector.scala 73:12]
    end else if (status == 8'h1) begin // @[Optimal_Weight_Vector.scala 75:26]
      status <= _status_T_1; // @[Optimal_Weight_Vector.scala 80:14]
    end else begin
      status <= _GEN_52;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  matrix_R_Comp_0_re = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  matrix_R_Comp_0_im = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  matrix_R_Comp_1_re = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  matrix_R_Comp_1_im = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  matrix_R_Comp_2_re = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  matrix_R_Comp_2_im = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  matrix_R_Comp_3_re = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  matrix_R_Comp_3_im = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  matrix_R_Comp_4_re = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  matrix_R_Comp_4_im = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  matrix_R_Comp_5_re = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  matrix_R_Comp_5_im = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  matrix_R_Comp_6_re = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  matrix_R_Comp_6_im = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  matrix_R_Comp_7_re = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  matrix_R_Comp_7_im = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  matrix_R_Comp_8_re = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  matrix_R_Comp_8_im = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  matrix_R_Comp_9_re = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  matrix_R_Comp_9_im = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  matrix_R_Comp_10_re = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  matrix_R_Comp_10_im = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  matrix_R_Comp_11_re = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  matrix_R_Comp_11_im = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  matrix_R_Comp_12_re = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  matrix_R_Comp_12_im = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  matrix_R_Comp_13_re = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  matrix_R_Comp_13_im = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  matrix_R_Comp_14_re = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  matrix_R_Comp_14_im = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  matrix_R_Comp_15_re = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  matrix_R_Comp_15_im = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  matrix_S_Comp_0_re = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  matrix_S_Comp_0_im = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  matrix_S_Comp_1_re = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  matrix_S_Comp_1_im = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  matrix_S_Comp_2_re = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  matrix_S_Comp_2_im = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  matrix_S_Comp_3_re = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  matrix_S_Comp_3_im = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  u_re = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  u_im = _RAND_41[63:0];
  _RAND_42 = {1{`RANDOM}};
  status = _RAND_42[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module matrix_conjugate_1(
  input  [63:0] io_matrixIn_0_re,
  input  [63:0] io_matrixIn_0_im,
  input  [63:0] io_matrixIn_4_re,
  input  [63:0] io_matrixIn_4_im,
  input  [63:0] io_matrixIn_5_re,
  input  [63:0] io_matrixIn_5_im,
  input  [63:0] io_matrixIn_8_re,
  input  [63:0] io_matrixIn_8_im,
  input  [63:0] io_matrixIn_9_re,
  input  [63:0] io_matrixIn_9_im,
  input  [63:0] io_matrixIn_10_re,
  input  [63:0] io_matrixIn_10_im,
  input  [63:0] io_matrixIn_12_re,
  input  [63:0] io_matrixIn_12_im,
  input  [63:0] io_matrixIn_13_re,
  input  [63:0] io_matrixIn_13_im,
  input  [63:0] io_matrixIn_14_re,
  input  [63:0] io_matrixIn_14_im,
  input  [63:0] io_matrixIn_15_re,
  input  [63:0] io_matrixIn_15_im,
  output [63:0] io_matrixOut_0_re,
  output [63:0] io_matrixOut_0_im,
  output [63:0] io_matrixOut_4_re,
  output [63:0] io_matrixOut_4_im,
  output [63:0] io_matrixOut_5_re,
  output [63:0] io_matrixOut_5_im,
  output [63:0] io_matrixOut_8_re,
  output [63:0] io_matrixOut_8_im,
  output [63:0] io_matrixOut_9_re,
  output [63:0] io_matrixOut_9_im,
  output [63:0] io_matrixOut_10_re,
  output [63:0] io_matrixOut_10_im,
  output [63:0] io_matrixOut_12_re,
  output [63:0] io_matrixOut_12_im,
  output [63:0] io_matrixOut_13_re,
  output [63:0] io_matrixOut_13_im,
  output [63:0] io_matrixOut_14_re,
  output [63:0] io_matrixOut_14_im,
  output [63:0] io_matrixOut_15_re,
  output [63:0] io_matrixOut_15_im
);
  assign io_matrixOut_0_re = io_matrixIn_0_re; // @[Matrix_Conjugate.scala 22:34]
  assign io_matrixOut_0_im = 64'sh0 - $signed(io_matrixIn_0_im); // @[Matrix_Conjugate.scala 23:37]
  assign io_matrixOut_4_re = io_matrixIn_4_re; // @[Matrix_Conjugate.scala 22:34]
  assign io_matrixOut_4_im = 64'sh0 - $signed(io_matrixIn_4_im); // @[Matrix_Conjugate.scala 23:37]
  assign io_matrixOut_5_re = io_matrixIn_5_re; // @[Matrix_Conjugate.scala 22:34]
  assign io_matrixOut_5_im = 64'sh0 - $signed(io_matrixIn_5_im); // @[Matrix_Conjugate.scala 23:37]
  assign io_matrixOut_8_re = io_matrixIn_8_re; // @[Matrix_Conjugate.scala 22:34]
  assign io_matrixOut_8_im = 64'sh0 - $signed(io_matrixIn_8_im); // @[Matrix_Conjugate.scala 23:37]
  assign io_matrixOut_9_re = io_matrixIn_9_re; // @[Matrix_Conjugate.scala 22:34]
  assign io_matrixOut_9_im = 64'sh0 - $signed(io_matrixIn_9_im); // @[Matrix_Conjugate.scala 23:37]
  assign io_matrixOut_10_re = io_matrixIn_10_re; // @[Matrix_Conjugate.scala 22:34]
  assign io_matrixOut_10_im = 64'sh0 - $signed(io_matrixIn_10_im); // @[Matrix_Conjugate.scala 23:37]
  assign io_matrixOut_12_re = io_matrixIn_12_re; // @[Matrix_Conjugate.scala 22:34]
  assign io_matrixOut_12_im = 64'sh0 - $signed(io_matrixIn_12_im); // @[Matrix_Conjugate.scala 23:37]
  assign io_matrixOut_13_re = io_matrixIn_13_re; // @[Matrix_Conjugate.scala 22:34]
  assign io_matrixOut_13_im = 64'sh0 - $signed(io_matrixIn_13_im); // @[Matrix_Conjugate.scala 23:37]
  assign io_matrixOut_14_re = io_matrixIn_14_re; // @[Matrix_Conjugate.scala 22:34]
  assign io_matrixOut_14_im = 64'sh0 - $signed(io_matrixIn_14_im); // @[Matrix_Conjugate.scala 23:37]
  assign io_matrixOut_15_re = io_matrixIn_15_re; // @[Matrix_Conjugate.scala 22:34]
  assign io_matrixOut_15_im = 64'sh0 - $signed(io_matrixIn_15_im); // @[Matrix_Conjugate.scala 23:37]
endmodule
module matrix_transpose_1(
  input  [63:0] io_matrixIn_0_re,
  input  [63:0] io_matrixIn_0_im,
  input  [63:0] io_matrixIn_4_re,
  input  [63:0] io_matrixIn_4_im,
  input  [63:0] io_matrixIn_5_re,
  input  [63:0] io_matrixIn_5_im,
  input  [63:0] io_matrixIn_8_re,
  input  [63:0] io_matrixIn_8_im,
  input  [63:0] io_matrixIn_9_re,
  input  [63:0] io_matrixIn_9_im,
  input  [63:0] io_matrixIn_10_re,
  input  [63:0] io_matrixIn_10_im,
  input  [63:0] io_matrixIn_12_re,
  input  [63:0] io_matrixIn_12_im,
  input  [63:0] io_matrixIn_13_re,
  input  [63:0] io_matrixIn_13_im,
  input  [63:0] io_matrixIn_14_re,
  input  [63:0] io_matrixIn_14_im,
  input  [63:0] io_matrixIn_15_re,
  input  [63:0] io_matrixIn_15_im,
  output [63:0] io_matrixOut_0_re,
  output [63:0] io_matrixOut_0_im,
  output [63:0] io_matrixOut_1_re,
  output [63:0] io_matrixOut_1_im,
  output [63:0] io_matrixOut_2_re,
  output [63:0] io_matrixOut_2_im,
  output [63:0] io_matrixOut_3_re,
  output [63:0] io_matrixOut_3_im,
  output [63:0] io_matrixOut_5_re,
  output [63:0] io_matrixOut_5_im,
  output [63:0] io_matrixOut_6_re,
  output [63:0] io_matrixOut_6_im,
  output [63:0] io_matrixOut_7_re,
  output [63:0] io_matrixOut_7_im,
  output [63:0] io_matrixOut_10_re,
  output [63:0] io_matrixOut_10_im,
  output [63:0] io_matrixOut_11_re,
  output [63:0] io_matrixOut_11_im,
  output [63:0] io_matrixOut_15_re,
  output [63:0] io_matrixOut_15_im
);
  assign io_matrixOut_0_re = io_matrixIn_0_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_0_im = io_matrixIn_0_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_1_re = io_matrixIn_4_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_1_im = io_matrixIn_4_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_2_re = io_matrixIn_8_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_2_im = io_matrixIn_8_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_3_re = io_matrixIn_12_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_3_im = io_matrixIn_12_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_5_re = io_matrixIn_5_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_5_im = io_matrixIn_5_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_6_re = io_matrixIn_9_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_6_im = io_matrixIn_9_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_7_re = io_matrixIn_13_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_7_im = io_matrixIn_13_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_10_re = io_matrixIn_10_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_10_im = io_matrixIn_10_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_11_re = io_matrixIn_14_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_11_im = io_matrixIn_14_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_15_re = io_matrixIn_15_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_15_im = io_matrixIn_15_im; // @[Matrix_Transpose.scala 22:31]
endmodule
module matirx_conjugate_transpose_1(
  input  [63:0] io_matrixIn_0_re,
  input  [63:0] io_matrixIn_0_im,
  input  [63:0] io_matrixIn_4_re,
  input  [63:0] io_matrixIn_4_im,
  input  [63:0] io_matrixIn_5_re,
  input  [63:0] io_matrixIn_5_im,
  input  [63:0] io_matrixIn_8_re,
  input  [63:0] io_matrixIn_8_im,
  input  [63:0] io_matrixIn_9_re,
  input  [63:0] io_matrixIn_9_im,
  input  [63:0] io_matrixIn_10_re,
  input  [63:0] io_matrixIn_10_im,
  input  [63:0] io_matrixIn_12_re,
  input  [63:0] io_matrixIn_12_im,
  input  [63:0] io_matrixIn_13_re,
  input  [63:0] io_matrixIn_13_im,
  input  [63:0] io_matrixIn_14_re,
  input  [63:0] io_matrixIn_14_im,
  input  [63:0] io_matrixIn_15_re,
  input  [63:0] io_matrixIn_15_im,
  output [63:0] io_matrixOut_0_re,
  output [63:0] io_matrixOut_0_im,
  output [63:0] io_matrixOut_1_re,
  output [63:0] io_matrixOut_1_im,
  output [63:0] io_matrixOut_2_re,
  output [63:0] io_matrixOut_2_im,
  output [63:0] io_matrixOut_3_re,
  output [63:0] io_matrixOut_3_im,
  output [63:0] io_matrixOut_5_re,
  output [63:0] io_matrixOut_5_im,
  output [63:0] io_matrixOut_6_re,
  output [63:0] io_matrixOut_6_im,
  output [63:0] io_matrixOut_7_re,
  output [63:0] io_matrixOut_7_im,
  output [63:0] io_matrixOut_10_re,
  output [63:0] io_matrixOut_10_im,
  output [63:0] io_matrixOut_11_re,
  output [63:0] io_matrixOut_11_im,
  output [63:0] io_matrixOut_15_re,
  output [63:0] io_matrixOut_15_im
);
  wire [63:0] unit_io_matrixIn_0_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_0_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_4_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_4_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_5_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_5_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_8_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_8_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_9_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_9_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_10_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_10_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_12_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_12_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_13_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_13_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_14_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_14_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_15_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixIn_15_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_0_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_0_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_4_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_4_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_5_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_5_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_8_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_8_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_9_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_9_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_10_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_10_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_12_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_12_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_13_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_13_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_14_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_14_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_15_re; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_io_matrixOut_15_im; // @[Matrix_Conjugate.scala 37:22]
  wire [63:0] unit_1_io_matrixIn_0_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_0_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_4_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_4_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_5_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_5_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_8_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_8_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_9_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_9_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_10_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_10_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_12_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_12_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_13_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_13_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_14_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_14_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_15_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixIn_15_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_0_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_0_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_1_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_1_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_2_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_2_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_3_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_3_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_5_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_5_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_6_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_6_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_7_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_7_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_10_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_10_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_11_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_11_im; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_15_re; // @[Matrix_Transpose.scala 36:22]
  wire [63:0] unit_1_io_matrixOut_15_im; // @[Matrix_Transpose.scala 36:22]
  matrix_conjugate_1 unit ( // @[Matrix_Conjugate.scala 37:22]
    .io_matrixIn_0_re(unit_io_matrixIn_0_re),
    .io_matrixIn_0_im(unit_io_matrixIn_0_im),
    .io_matrixIn_4_re(unit_io_matrixIn_4_re),
    .io_matrixIn_4_im(unit_io_matrixIn_4_im),
    .io_matrixIn_5_re(unit_io_matrixIn_5_re),
    .io_matrixIn_5_im(unit_io_matrixIn_5_im),
    .io_matrixIn_8_re(unit_io_matrixIn_8_re),
    .io_matrixIn_8_im(unit_io_matrixIn_8_im),
    .io_matrixIn_9_re(unit_io_matrixIn_9_re),
    .io_matrixIn_9_im(unit_io_matrixIn_9_im),
    .io_matrixIn_10_re(unit_io_matrixIn_10_re),
    .io_matrixIn_10_im(unit_io_matrixIn_10_im),
    .io_matrixIn_12_re(unit_io_matrixIn_12_re),
    .io_matrixIn_12_im(unit_io_matrixIn_12_im),
    .io_matrixIn_13_re(unit_io_matrixIn_13_re),
    .io_matrixIn_13_im(unit_io_matrixIn_13_im),
    .io_matrixIn_14_re(unit_io_matrixIn_14_re),
    .io_matrixIn_14_im(unit_io_matrixIn_14_im),
    .io_matrixIn_15_re(unit_io_matrixIn_15_re),
    .io_matrixIn_15_im(unit_io_matrixIn_15_im),
    .io_matrixOut_0_re(unit_io_matrixOut_0_re),
    .io_matrixOut_0_im(unit_io_matrixOut_0_im),
    .io_matrixOut_4_re(unit_io_matrixOut_4_re),
    .io_matrixOut_4_im(unit_io_matrixOut_4_im),
    .io_matrixOut_5_re(unit_io_matrixOut_5_re),
    .io_matrixOut_5_im(unit_io_matrixOut_5_im),
    .io_matrixOut_8_re(unit_io_matrixOut_8_re),
    .io_matrixOut_8_im(unit_io_matrixOut_8_im),
    .io_matrixOut_9_re(unit_io_matrixOut_9_re),
    .io_matrixOut_9_im(unit_io_matrixOut_9_im),
    .io_matrixOut_10_re(unit_io_matrixOut_10_re),
    .io_matrixOut_10_im(unit_io_matrixOut_10_im),
    .io_matrixOut_12_re(unit_io_matrixOut_12_re),
    .io_matrixOut_12_im(unit_io_matrixOut_12_im),
    .io_matrixOut_13_re(unit_io_matrixOut_13_re),
    .io_matrixOut_13_im(unit_io_matrixOut_13_im),
    .io_matrixOut_14_re(unit_io_matrixOut_14_re),
    .io_matrixOut_14_im(unit_io_matrixOut_14_im),
    .io_matrixOut_15_re(unit_io_matrixOut_15_re),
    .io_matrixOut_15_im(unit_io_matrixOut_15_im)
  );
  matrix_transpose_1 unit_1 ( // @[Matrix_Transpose.scala 36:22]
    .io_matrixIn_0_re(unit_1_io_matrixIn_0_re),
    .io_matrixIn_0_im(unit_1_io_matrixIn_0_im),
    .io_matrixIn_4_re(unit_1_io_matrixIn_4_re),
    .io_matrixIn_4_im(unit_1_io_matrixIn_4_im),
    .io_matrixIn_5_re(unit_1_io_matrixIn_5_re),
    .io_matrixIn_5_im(unit_1_io_matrixIn_5_im),
    .io_matrixIn_8_re(unit_1_io_matrixIn_8_re),
    .io_matrixIn_8_im(unit_1_io_matrixIn_8_im),
    .io_matrixIn_9_re(unit_1_io_matrixIn_9_re),
    .io_matrixIn_9_im(unit_1_io_matrixIn_9_im),
    .io_matrixIn_10_re(unit_1_io_matrixIn_10_re),
    .io_matrixIn_10_im(unit_1_io_matrixIn_10_im),
    .io_matrixIn_12_re(unit_1_io_matrixIn_12_re),
    .io_matrixIn_12_im(unit_1_io_matrixIn_12_im),
    .io_matrixIn_13_re(unit_1_io_matrixIn_13_re),
    .io_matrixIn_13_im(unit_1_io_matrixIn_13_im),
    .io_matrixIn_14_re(unit_1_io_matrixIn_14_re),
    .io_matrixIn_14_im(unit_1_io_matrixIn_14_im),
    .io_matrixIn_15_re(unit_1_io_matrixIn_15_re),
    .io_matrixIn_15_im(unit_1_io_matrixIn_15_im),
    .io_matrixOut_0_re(unit_1_io_matrixOut_0_re),
    .io_matrixOut_0_im(unit_1_io_matrixOut_0_im),
    .io_matrixOut_1_re(unit_1_io_matrixOut_1_re),
    .io_matrixOut_1_im(unit_1_io_matrixOut_1_im),
    .io_matrixOut_2_re(unit_1_io_matrixOut_2_re),
    .io_matrixOut_2_im(unit_1_io_matrixOut_2_im),
    .io_matrixOut_3_re(unit_1_io_matrixOut_3_re),
    .io_matrixOut_3_im(unit_1_io_matrixOut_3_im),
    .io_matrixOut_5_re(unit_1_io_matrixOut_5_re),
    .io_matrixOut_5_im(unit_1_io_matrixOut_5_im),
    .io_matrixOut_6_re(unit_1_io_matrixOut_6_re),
    .io_matrixOut_6_im(unit_1_io_matrixOut_6_im),
    .io_matrixOut_7_re(unit_1_io_matrixOut_7_re),
    .io_matrixOut_7_im(unit_1_io_matrixOut_7_im),
    .io_matrixOut_10_re(unit_1_io_matrixOut_10_re),
    .io_matrixOut_10_im(unit_1_io_matrixOut_10_im),
    .io_matrixOut_11_re(unit_1_io_matrixOut_11_re),
    .io_matrixOut_11_im(unit_1_io_matrixOut_11_im),
    .io_matrixOut_15_re(unit_1_io_matrixOut_15_re),
    .io_matrixOut_15_im(unit_1_io_matrixOut_15_im)
  );
  assign io_matrixOut_0_re = unit_1_io_matrixOut_0_re; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_0_im = unit_1_io_matrixOut_0_im; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_1_re = unit_1_io_matrixOut_1_re; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_1_im = unit_1_io_matrixOut_1_im; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_2_re = unit_1_io_matrixOut_2_re; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_2_im = unit_1_io_matrixOut_2_im; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_3_re = unit_1_io_matrixOut_3_re; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_3_im = unit_1_io_matrixOut_3_im; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_5_re = unit_1_io_matrixOut_5_re; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_5_im = unit_1_io_matrixOut_5_im; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_6_re = unit_1_io_matrixOut_6_re; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_6_im = unit_1_io_matrixOut_6_im; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_7_re = unit_1_io_matrixOut_7_re; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_7_im = unit_1_io_matrixOut_7_im; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_10_re = unit_1_io_matrixOut_10_re; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_10_im = unit_1_io_matrixOut_10_im; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_11_re = unit_1_io_matrixOut_11_re; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_11_im = unit_1_io_matrixOut_11_im; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_15_re = unit_1_io_matrixOut_15_re; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign io_matrixOut_15_im = unit_1_io_matrixOut_15_im; // @[Matirx_Conjugate_Transpose.scala 20:16]
  assign unit_io_matrixIn_0_re = io_matrixIn_0_re; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_0_im = io_matrixIn_0_im; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_4_re = io_matrixIn_4_re; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_4_im = io_matrixIn_4_im; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_5_re = io_matrixIn_5_re; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_5_im = io_matrixIn_5_im; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_8_re = io_matrixIn_8_re; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_8_im = io_matrixIn_8_im; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_9_re = io_matrixIn_9_re; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_9_im = io_matrixIn_9_im; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_10_re = io_matrixIn_10_re; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_10_im = io_matrixIn_10_im; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_12_re = io_matrixIn_12_re; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_12_im = io_matrixIn_12_im; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_13_re = io_matrixIn_13_re; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_13_im = io_matrixIn_13_im; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_14_re = io_matrixIn_14_re; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_14_im = io_matrixIn_14_im; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_15_re = io_matrixIn_15_re; // @[Matrix_Conjugate.scala 38:22]
  assign unit_io_matrixIn_15_im = io_matrixIn_15_im; // @[Matrix_Conjugate.scala 38:22]
  assign unit_1_io_matrixIn_0_re = unit_io_matrixOut_0_re; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_0_im = unit_io_matrixOut_0_im; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_4_re = unit_io_matrixOut_4_re; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_4_im = unit_io_matrixOut_4_im; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_5_re = unit_io_matrixOut_5_re; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_5_im = unit_io_matrixOut_5_im; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_8_re = unit_io_matrixOut_8_re; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_8_im = unit_io_matrixOut_8_im; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_9_re = unit_io_matrixOut_9_re; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_9_im = unit_io_matrixOut_9_im; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_10_re = unit_io_matrixOut_10_re; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_10_im = unit_io_matrixOut_10_im; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_12_re = unit_io_matrixOut_12_re; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_12_im = unit_io_matrixOut_12_im; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_13_re = unit_io_matrixOut_13_re; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_13_im = unit_io_matrixOut_13_im; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_14_re = unit_io_matrixOut_14_re; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_14_im = unit_io_matrixOut_14_im; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_15_re = unit_io_matrixOut_15_re; // @[Matrix_Transpose.scala 37:22]
  assign unit_1_io_matrixIn_15_im = unit_io_matrixOut_15_im; // @[Matrix_Transpose.scala 37:22]
endmodule
module stap_main(
  input         clock,
  input         reset,
  input         io_reset,
  input         io_ready,
  input  [63:0] io_theta,
  input  [63:0] io_psi,
  input  [63:0] io_d,
  input  [63:0] io_lambda,
  input  [63:0] io_v,
  input  [63:0] io_T,
  input  [63:0] io_matrixIn_0_re,
  input  [63:0] io_matrixIn_0_im,
  input  [63:0] io_matrixIn_1_re,
  input  [63:0] io_matrixIn_1_im,
  input  [63:0] io_matrixIn_2_re,
  input  [63:0] io_matrixIn_2_im,
  input  [63:0] io_matrixIn_3_re,
  input  [63:0] io_matrixIn_3_im,
  input  [63:0] io_matrixIn_4_re,
  input  [63:0] io_matrixIn_4_im,
  input  [63:0] io_matrixIn_5_re,
  input  [63:0] io_matrixIn_5_im,
  input  [63:0] io_matrixIn_6_re,
  input  [63:0] io_matrixIn_6_im,
  input  [63:0] io_matrixIn_7_re,
  input  [63:0] io_matrixIn_7_im,
  output [63:0] io_matrixOut_0_re,
  output [63:0] io_matrixOut_0_im,
  output [63:0] io_matrixOut_1_re,
  output [63:0] io_matrixOut_1_im,
  output [63:0] io_matrixOut_2_re,
  output [63:0] io_matrixOut_2_im,
  output [63:0] io_matrixOut_3_re,
  output [63:0] io_matrixOut_3_im,
  output        io_valid,
  output [7:0]  io_debug_status,
  output        io_debug_valid_R_matirx_estimation,
  output        io_debug_valid_cholesky_v1,
  output        io_debug_valid_lower_triangular_matrix_inversion_complex_v1,
  output        io_debug_valid_matrix_mul_v1,
  output        io_debug_valid_optimal_weight_vector,
  output [63:0] io_debug_matrix_x_in_0_re,
  output [63:0] io_debug_matrix_x_in_0_im,
  output [63:0] io_debug_matrix_x_in_1_re,
  output [63:0] io_debug_matrix_x_in_1_im,
  output [63:0] io_debug_matrix_x_in_2_re,
  output [63:0] io_debug_matrix_x_in_2_im,
  output [63:0] io_debug_matrix_x_in_3_re,
  output [63:0] io_debug_matrix_x_in_3_im,
  output [63:0] io_debug_matrix_x_in_4_re,
  output [63:0] io_debug_matrix_x_in_4_im,
  output [63:0] io_debug_matrix_x_in_5_re,
  output [63:0] io_debug_matrix_x_in_5_im,
  output [63:0] io_debug_matrix_x_in_6_re,
  output [63:0] io_debug_matrix_x_in_6_im,
  output [63:0] io_debug_matrix_x_in_7_re,
  output [63:0] io_debug_matrix_x_in_7_im,
  output [63:0] io_debug_matrix_S_0_re,
  output [63:0] io_debug_matrix_S_0_im,
  output [63:0] io_debug_matrix_S_1_re,
  output [63:0] io_debug_matrix_S_1_im,
  output [63:0] io_debug_matrix_S_2_re,
  output [63:0] io_debug_matrix_S_2_im,
  output [63:0] io_debug_matrix_S_3_re,
  output [63:0] io_debug_matrix_S_3_im,
  output [63:0] io_debug_matrix_R_0_re,
  output [63:0] io_debug_matrix_R_0_im,
  output [63:0] io_debug_matrix_R_1_re,
  output [63:0] io_debug_matrix_R_1_im,
  output [63:0] io_debug_matrix_R_2_re,
  output [63:0] io_debug_matrix_R_2_im,
  output [63:0] io_debug_matrix_R_3_re,
  output [63:0] io_debug_matrix_R_3_im,
  output [63:0] io_debug_matrix_R_4_re,
  output [63:0] io_debug_matrix_R_4_im,
  output [63:0] io_debug_matrix_R_5_re,
  output [63:0] io_debug_matrix_R_5_im,
  output [63:0] io_debug_matrix_R_6_re,
  output [63:0] io_debug_matrix_R_6_im,
  output [63:0] io_debug_matrix_R_7_re,
  output [63:0] io_debug_matrix_R_7_im,
  output [63:0] io_debug_matrix_R_8_re,
  output [63:0] io_debug_matrix_R_8_im,
  output [63:0] io_debug_matrix_R_9_re,
  output [63:0] io_debug_matrix_R_9_im,
  output [63:0] io_debug_matrix_R_10_re,
  output [63:0] io_debug_matrix_R_10_im,
  output [63:0] io_debug_matrix_R_11_re,
  output [63:0] io_debug_matrix_R_11_im,
  output [63:0] io_debug_matrix_R_12_re,
  output [63:0] io_debug_matrix_R_12_im,
  output [63:0] io_debug_matrix_R_13_re,
  output [63:0] io_debug_matrix_R_13_im,
  output [63:0] io_debug_matrix_R_14_re,
  output [63:0] io_debug_matrix_R_14_im,
  output [63:0] io_debug_matrix_R_15_re,
  output [63:0] io_debug_matrix_R_15_im,
  output [63:0] io_debug_matrix_L_0_re,
  output [63:0] io_debug_matrix_L_0_im,
  output [63:0] io_debug_matrix_L_1_re,
  output [63:0] io_debug_matrix_L_1_im,
  output [63:0] io_debug_matrix_L_2_re,
  output [63:0] io_debug_matrix_L_2_im,
  output [63:0] io_debug_matrix_L_3_re,
  output [63:0] io_debug_matrix_L_3_im,
  output [63:0] io_debug_matrix_L_4_re,
  output [63:0] io_debug_matrix_L_4_im,
  output [63:0] io_debug_matrix_L_5_re,
  output [63:0] io_debug_matrix_L_5_im,
  output [63:0] io_debug_matrix_L_6_re,
  output [63:0] io_debug_matrix_L_6_im,
  output [63:0] io_debug_matrix_L_7_re,
  output [63:0] io_debug_matrix_L_7_im,
  output [63:0] io_debug_matrix_L_8_re,
  output [63:0] io_debug_matrix_L_8_im,
  output [63:0] io_debug_matrix_L_9_re,
  output [63:0] io_debug_matrix_L_9_im,
  output [63:0] io_debug_matrix_L_inv_0_re,
  output [63:0] io_debug_matrix_L_inv_0_im,
  output [63:0] io_debug_matrix_L_inv_1_re,
  output [63:0] io_debug_matrix_L_inv_1_im,
  output [63:0] io_debug_matrix_L_inv_2_re,
  output [63:0] io_debug_matrix_L_inv_2_im,
  output [63:0] io_debug_matrix_L_inv_3_re,
  output [63:0] io_debug_matrix_L_inv_3_im,
  output [63:0] io_debug_matrix_L_inv_4_re,
  output [63:0] io_debug_matrix_L_inv_4_im,
  output [63:0] io_debug_matrix_L_inv_5_re,
  output [63:0] io_debug_matrix_L_inv_5_im,
  output [63:0] io_debug_matrix_L_inv_6_re,
  output [63:0] io_debug_matrix_L_inv_6_im,
  output [63:0] io_debug_matrix_L_inv_7_re,
  output [63:0] io_debug_matrix_L_inv_7_im,
  output [63:0] io_debug_matrix_L_inv_8_re,
  output [63:0] io_debug_matrix_L_inv_8_im,
  output [63:0] io_debug_matrix_L_inv_9_re,
  output [63:0] io_debug_matrix_L_inv_9_im,
  output [63:0] io_debug_matrix_R_inv_0_re,
  output [63:0] io_debug_matrix_R_inv_0_im,
  output [63:0] io_debug_matrix_R_inv_1_re,
  output [63:0] io_debug_matrix_R_inv_1_im,
  output [63:0] io_debug_matrix_R_inv_2_re,
  output [63:0] io_debug_matrix_R_inv_2_im,
  output [63:0] io_debug_matrix_R_inv_3_re,
  output [63:0] io_debug_matrix_R_inv_3_im,
  output [63:0] io_debug_matrix_R_inv_4_re,
  output [63:0] io_debug_matrix_R_inv_4_im,
  output [63:0] io_debug_matrix_R_inv_5_re,
  output [63:0] io_debug_matrix_R_inv_5_im,
  output [63:0] io_debug_matrix_R_inv_6_re,
  output [63:0] io_debug_matrix_R_inv_6_im,
  output [63:0] io_debug_matrix_R_inv_7_re,
  output [63:0] io_debug_matrix_R_inv_7_im,
  output [63:0] io_debug_matrix_R_inv_8_re,
  output [63:0] io_debug_matrix_R_inv_8_im,
  output [63:0] io_debug_matrix_R_inv_9_re,
  output [63:0] io_debug_matrix_R_inv_9_im,
  output [63:0] io_debug_matrix_R_inv_10_re,
  output [63:0] io_debug_matrix_R_inv_10_im,
  output [63:0] io_debug_matrix_R_inv_11_re,
  output [63:0] io_debug_matrix_R_inv_11_im,
  output [63:0] io_debug_matrix_R_inv_12_re,
  output [63:0] io_debug_matrix_R_inv_12_im,
  output [63:0] io_debug_matrix_R_inv_13_re,
  output [63:0] io_debug_matrix_R_inv_13_im,
  output [63:0] io_debug_matrix_R_inv_14_re,
  output [63:0] io_debug_matrix_R_inv_14_im,
  output [63:0] io_debug_matrix_R_inv_15_re,
  output [63:0] io_debug_matrix_R_inv_15_im,
  output [63:0] io_debug_matrix_w_0_re,
  output [63:0] io_debug_matrix_w_0_im,
  output [63:0] io_debug_matrix_w_1_re,
  output [63:0] io_debug_matrix_w_1_im,
  output [63:0] io_debug_matrix_w_2_re,
  output [63:0] io_debug_matrix_w_2_im,
  output [63:0] io_debug_matrix_w_3_re,
  output [63:0] io_debug_matrix_w_3_im
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [31:0] _RAND_136;
`endif // RANDOMIZE_REG_INIT
  wire  space_time_steering_vector_unit_clock; // @[Stap_Main.scala 81:47]
  wire  space_time_steering_vector_unit_reset; // @[Stap_Main.scala 81:47]
  wire [63:0] space_time_steering_vector_unit_io_theta; // @[Stap_Main.scala 81:47]
  wire [63:0] space_time_steering_vector_unit_io_psi; // @[Stap_Main.scala 81:47]
  wire [63:0] space_time_steering_vector_unit_io_d; // @[Stap_Main.scala 81:47]
  wire [63:0] space_time_steering_vector_unit_io_lambda; // @[Stap_Main.scala 81:47]
  wire [63:0] space_time_steering_vector_unit_io_v; // @[Stap_Main.scala 81:47]
  wire [63:0] space_time_steering_vector_unit_io_T; // @[Stap_Main.scala 81:47]
  wire [63:0] space_time_steering_vector_unit_io_matrixOut_0_re; // @[Stap_Main.scala 81:47]
  wire [63:0] space_time_steering_vector_unit_io_matrixOut_0_im; // @[Stap_Main.scala 81:47]
  wire [63:0] space_time_steering_vector_unit_io_matrixOut_1_re; // @[Stap_Main.scala 81:47]
  wire [63:0] space_time_steering_vector_unit_io_matrixOut_1_im; // @[Stap_Main.scala 81:47]
  wire [63:0] space_time_steering_vector_unit_io_matrixOut_2_re; // @[Stap_Main.scala 81:47]
  wire [63:0] space_time_steering_vector_unit_io_matrixOut_2_im; // @[Stap_Main.scala 81:47]
  wire [63:0] space_time_steering_vector_unit_io_matrixOut_3_re; // @[Stap_Main.scala 81:47]
  wire [63:0] space_time_steering_vector_unit_io_matrixOut_3_im; // @[Stap_Main.scala 81:47]
  wire  R_matirx_estimation_clock; // @[Stap_Main.scala 91:56]
  wire  R_matirx_estimation_reset; // @[Stap_Main.scala 91:56]
  wire  R_matirx_estimation_io_reset; // @[Stap_Main.scala 91:56]
  wire  R_matirx_estimation_io_ready; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixIn_0_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixIn_0_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixIn_1_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixIn_1_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixIn_2_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixIn_2_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixIn_3_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixIn_3_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixIn_4_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixIn_4_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixIn_5_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixIn_5_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixIn_6_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixIn_6_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixIn_7_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixIn_7_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_0_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_0_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_1_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_1_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_2_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_2_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_3_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_3_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_4_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_4_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_5_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_5_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_6_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_6_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_7_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_7_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_8_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_8_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_9_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_9_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_10_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_10_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_11_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_11_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_12_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_12_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_13_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_13_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_14_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_14_im; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_15_re; // @[Stap_Main.scala 91:56]
  wire [63:0] R_matirx_estimation_io_matrixOut_15_im; // @[Stap_Main.scala 91:56]
  wire  R_matirx_estimation_io_valid; // @[Stap_Main.scala 91:56]
  wire  cholesky_v1_clock; // @[Stap_Main.scala 92:40]
  wire  cholesky_v1_reset; // @[Stap_Main.scala 92:40]
  wire  cholesky_v1_io_reset; // @[Stap_Main.scala 92:40]
  wire  cholesky_v1_io_ready; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_0_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_0_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_1_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_1_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_2_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_2_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_3_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_3_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_4_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_4_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_5_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_5_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_6_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_6_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_7_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_7_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_8_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_8_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_9_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_9_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_10_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_10_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_11_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_11_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_12_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_12_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_13_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_13_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_14_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_14_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_15_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixIn_15_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_0_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_0_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_1_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_1_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_2_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_2_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_3_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_3_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_4_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_4_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_5_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_5_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_6_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_6_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_7_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_7_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_8_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_8_im; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_9_re; // @[Stap_Main.scala 92:40]
  wire [63:0] cholesky_v1_io_matrixOut_9_im; // @[Stap_Main.scala 92:40]
  wire  cholesky_v1_io_valid; // @[Stap_Main.scala 92:40]
  wire  lower_triangular_matrix_inversion_complex_v1_clock; // @[Stap_Main.scala 93:60]
  wire  lower_triangular_matrix_inversion_complex_v1_reset; // @[Stap_Main.scala 93:60]
  wire  lower_triangular_matrix_inversion_complex_v1_io_reset; // @[Stap_Main.scala 93:60]
  wire  lower_triangular_matrix_inversion_complex_v1_io_ready; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_0_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_0_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_1_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_1_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_2_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_2_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_3_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_3_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_4_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_4_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_5_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_5_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_6_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_6_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_7_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_7_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_8_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_8_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_9_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixIn_9_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_0_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_0_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_1_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_1_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_2_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_2_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_3_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_3_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_4_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_4_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_5_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_5_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_6_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_6_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_7_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_7_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_8_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_8_im; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_9_re; // @[Stap_Main.scala 93:60]
  wire [63:0] lower_triangular_matrix_inversion_complex_v1_io_matrixOut_9_im; // @[Stap_Main.scala 93:60]
  wire  lower_triangular_matrix_inversion_complex_v1_io_valid; // @[Stap_Main.scala 93:60]
  wire  matrix_mul_v1_clock; // @[Stap_Main.scala 94:44]
  wire  matrix_mul_v1_io_reset; // @[Stap_Main.scala 94:44]
  wire  matrix_mul_v1_io_ready; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_0_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_0_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_1_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_1_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_2_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_2_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_3_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_3_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_5_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_5_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_6_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_6_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_7_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_7_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_10_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_10_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_11_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_11_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_15_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixA_15_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_0_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_0_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_4_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_4_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_5_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_5_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_8_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_8_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_9_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_9_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_10_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_10_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_12_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_12_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_13_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_13_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_14_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_14_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_15_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixB_15_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_0_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_0_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_1_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_1_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_2_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_2_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_3_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_3_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_4_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_4_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_5_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_5_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_6_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_6_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_7_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_7_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_8_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_8_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_9_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_9_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_10_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_10_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_11_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_11_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_12_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_12_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_13_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_13_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_14_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_14_im; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_15_re; // @[Stap_Main.scala 94:44]
  wire [63:0] matrix_mul_v1_io_matrixC_15_im; // @[Stap_Main.scala 94:44]
  wire  matrix_mul_v1_io_valid; // @[Stap_Main.scala 94:44]
  wire  optimal_weight_vector_clock; // @[Stap_Main.scala 95:60]
  wire  optimal_weight_vector_reset; // @[Stap_Main.scala 95:60]
  wire  optimal_weight_vector_io_reset; // @[Stap_Main.scala 95:60]
  wire  optimal_weight_vector_io_ready; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixS_0_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixS_0_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixS_1_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixS_1_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixS_2_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixS_2_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixS_3_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixS_3_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_0_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_0_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_1_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_1_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_2_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_2_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_3_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_3_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_4_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_4_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_5_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_5_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_6_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_6_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_7_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_7_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_8_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_8_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_9_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_9_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_10_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_10_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_11_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_11_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_12_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_12_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_13_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_13_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_14_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_14_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_15_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixR_Inv_15_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixOut_0_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixOut_0_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixOut_1_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixOut_1_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixOut_2_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixOut_2_im; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixOut_3_re; // @[Stap_Main.scala 95:60]
  wire [63:0] optimal_weight_vector_io_matrixOut_3_im; // @[Stap_Main.scala 95:60]
  wire  optimal_weight_vector_io_valid; // @[Stap_Main.scala 95:60]
  wire [63:0] unit_io_matrixIn_0_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_0_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_4_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_4_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_5_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_5_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_8_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_8_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_9_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_9_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_10_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_10_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_12_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_12_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_13_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_13_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_14_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_14_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_15_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixIn_15_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_0_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_0_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_1_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_1_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_2_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_2_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_3_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_3_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_5_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_5_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_6_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_6_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_7_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_7_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_10_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_10_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_11_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_11_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_15_re; // @[Matirx_Conjugate_Transpose.scala 32:22]
  wire [63:0] unit_io_matrixOut_15_im; // @[Matirx_Conjugate_Transpose.scala 32:22]
  reg [63:0] matrix_x_in_0_re; // @[Stap_Main.scala 59:38]
  reg [63:0] matrix_x_in_0_im; // @[Stap_Main.scala 59:38]
  reg [63:0] matrix_x_in_1_re; // @[Stap_Main.scala 59:38]
  reg [63:0] matrix_x_in_1_im; // @[Stap_Main.scala 59:38]
  reg [63:0] matrix_x_in_2_re; // @[Stap_Main.scala 59:38]
  reg [63:0] matrix_x_in_2_im; // @[Stap_Main.scala 59:38]
  reg [63:0] matrix_x_in_3_re; // @[Stap_Main.scala 59:38]
  reg [63:0] matrix_x_in_3_im; // @[Stap_Main.scala 59:38]
  reg [63:0] matrix_x_in_4_re; // @[Stap_Main.scala 59:38]
  reg [63:0] matrix_x_in_4_im; // @[Stap_Main.scala 59:38]
  reg [63:0] matrix_x_in_5_re; // @[Stap_Main.scala 59:38]
  reg [63:0] matrix_x_in_5_im; // @[Stap_Main.scala 59:38]
  reg [63:0] matrix_x_in_6_re; // @[Stap_Main.scala 59:38]
  reg [63:0] matrix_x_in_6_im; // @[Stap_Main.scala 59:38]
  reg [63:0] matrix_x_in_7_re; // @[Stap_Main.scala 59:38]
  reg [63:0] matrix_x_in_7_im; // @[Stap_Main.scala 59:38]
  reg [63:0] matrix_S_0_re; // @[Stap_Main.scala 60:35]
  reg [63:0] matrix_S_0_im; // @[Stap_Main.scala 60:35]
  reg [63:0] matrix_S_1_re; // @[Stap_Main.scala 60:35]
  reg [63:0] matrix_S_1_im; // @[Stap_Main.scala 60:35]
  reg [63:0] matrix_S_2_re; // @[Stap_Main.scala 60:35]
  reg [63:0] matrix_S_2_im; // @[Stap_Main.scala 60:35]
  reg [63:0] matrix_S_3_re; // @[Stap_Main.scala 60:35]
  reg [63:0] matrix_S_3_im; // @[Stap_Main.scala 60:35]
  reg [63:0] matrix_R_0_re; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_0_im; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_1_re; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_1_im; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_2_re; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_2_im; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_3_re; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_3_im; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_4_re; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_4_im; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_5_re; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_5_im; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_6_re; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_6_im; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_7_re; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_7_im; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_8_re; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_8_im; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_9_re; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_9_im; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_10_re; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_10_im; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_11_re; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_11_im; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_12_re; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_12_im; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_13_re; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_13_im; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_14_re; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_14_im; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_15_re; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_R_15_im; // @[Stap_Main.scala 61:35]
  reg [63:0] matrix_L_0_re; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_0_im; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_1_re; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_1_im; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_2_re; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_2_im; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_3_re; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_3_im; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_4_re; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_4_im; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_5_re; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_5_im; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_6_re; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_6_im; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_7_re; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_7_im; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_8_re; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_8_im; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_9_re; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_9_im; // @[Stap_Main.scala 62:35]
  reg [63:0] matrix_L_inv_0_re; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_0_im; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_1_re; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_1_im; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_2_re; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_2_im; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_3_re; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_3_im; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_4_re; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_4_im; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_5_re; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_5_im; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_6_re; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_6_im; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_7_re; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_7_im; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_8_re; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_8_im; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_9_re; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_L_inv_9_im; // @[Stap_Main.scala 63:39]
  reg [63:0] matrix_R_inv_0_re; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_0_im; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_1_re; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_1_im; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_2_re; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_2_im; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_3_re; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_3_im; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_4_re; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_4_im; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_5_re; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_5_im; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_6_re; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_6_im; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_7_re; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_7_im; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_8_re; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_8_im; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_9_re; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_9_im; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_10_re; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_10_im; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_11_re; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_11_im; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_12_re; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_12_im; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_13_re; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_13_im; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_14_re; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_14_im; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_15_re; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_R_inv_15_im; // @[Stap_Main.scala 64:39]
  reg [63:0] matrix_w_0_re; // @[Stap_Main.scala 65:35]
  reg [63:0] matrix_w_0_im; // @[Stap_Main.scala 65:35]
  reg [63:0] matrix_w_1_re; // @[Stap_Main.scala 65:35]
  reg [63:0] matrix_w_1_im; // @[Stap_Main.scala 65:35]
  reg [63:0] matrix_w_2_re; // @[Stap_Main.scala 65:35]
  reg [63:0] matrix_w_2_im; // @[Stap_Main.scala 65:35]
  reg [63:0] matrix_w_3_re; // @[Stap_Main.scala 65:35]
  reg [63:0] matrix_w_3_im; // @[Stap_Main.scala 65:35]
  reg [7:0] status; // @[Stap_Main.scala 66:29]
  wire [7:0] _status_T_1 = status + 8'h1; // @[Stap_Main.scala 146:24]
  wire [63:0] _GEN_0 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_0_im) : $signed(
    matrix_R_0_im); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_1 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_0_re) : $signed(
    matrix_R_0_re); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_2 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_1_im) : $signed(
    matrix_R_1_im); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_3 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_1_re) : $signed(
    matrix_R_1_re); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_4 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_2_im) : $signed(
    matrix_R_2_im); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_5 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_2_re) : $signed(
    matrix_R_2_re); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_6 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_3_im) : $signed(
    matrix_R_3_im); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_7 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_3_re) : $signed(
    matrix_R_3_re); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_8 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_4_im) : $signed(
    matrix_R_4_im); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_9 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_4_re) : $signed(
    matrix_R_4_re); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_10 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_5_im) : $signed(
    matrix_R_5_im); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_11 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_5_re) : $signed(
    matrix_R_5_re); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_12 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_6_im) : $signed(
    matrix_R_6_im); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_13 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_6_re) : $signed(
    matrix_R_6_re); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_14 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_7_im) : $signed(
    matrix_R_7_im); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_15 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_7_re) : $signed(
    matrix_R_7_re); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_16 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_8_im) : $signed(
    matrix_R_8_im); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_17 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_8_re) : $signed(
    matrix_R_8_re); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_18 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_9_im) : $signed(
    matrix_R_9_im); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_19 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_9_re) : $signed(
    matrix_R_9_re); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_20 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_10_im) : $signed(
    matrix_R_10_im); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_21 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_10_re) : $signed(
    matrix_R_10_re); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_22 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_11_im) : $signed(
    matrix_R_11_im); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_23 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_11_re) : $signed(
    matrix_R_11_re); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_24 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_12_im) : $signed(
    matrix_R_12_im); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_25 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_12_re) : $signed(
    matrix_R_12_re); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_26 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_13_im) : $signed(
    matrix_R_13_im); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_27 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_13_re) : $signed(
    matrix_R_13_re); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_28 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_14_im) : $signed(
    matrix_R_14_im); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_29 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_14_re) : $signed(
    matrix_R_14_re); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_30 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_15_im) : $signed(
    matrix_R_15_im); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [63:0] _GEN_31 = R_matirx_estimation_io_valid ? $signed(R_matirx_estimation_io_matrixOut_15_re) : $signed(
    matrix_R_15_re); // @[Stap_Main.scala 150:42 151:18 61:35]
  wire [7:0] _GEN_32 = R_matirx_estimation_io_valid ? _status_T_1 : status; // @[Stap_Main.scala 150:42 152:16 66:29]
  wire [63:0] _GEN_33 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_0_im) : $signed(matrix_L_0_im); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_34 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_0_re) : $signed(matrix_L_0_re); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_35 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_1_im) : $signed(matrix_L_1_im); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_36 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_1_re) : $signed(matrix_L_1_re); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_37 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_2_im) : $signed(matrix_L_2_im); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_38 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_2_re) : $signed(matrix_L_2_re); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_39 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_3_im) : $signed(matrix_L_3_im); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_40 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_3_re) : $signed(matrix_L_3_re); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_41 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_4_im) : $signed(matrix_L_4_im); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_42 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_4_re) : $signed(matrix_L_4_re); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_43 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_5_im) : $signed(matrix_L_5_im); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_44 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_5_re) : $signed(matrix_L_5_re); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_45 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_6_im) : $signed(matrix_L_6_im); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_46 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_6_re) : $signed(matrix_L_6_re); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_47 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_7_im) : $signed(matrix_L_7_im); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_48 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_7_re) : $signed(matrix_L_7_re); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_49 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_8_im) : $signed(matrix_L_8_im); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_50 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_8_re) : $signed(matrix_L_8_re); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_51 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_9_im) : $signed(matrix_L_9_im); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [63:0] _GEN_52 = cholesky_v1_io_valid ? $signed(cholesky_v1_io_matrixOut_9_re) : $signed(matrix_L_9_re); // @[Stap_Main.scala 162:34 163:18 62:35]
  wire [7:0] _GEN_53 = cholesky_v1_io_valid ? _status_T_1 : status; // @[Stap_Main.scala 162:34 164:16 66:29]
  wire [63:0] _GEN_54 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_0_im) : $signed(matrix_L_inv_0_im); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_55 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_0_re) : $signed(matrix_L_inv_0_re); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_56 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_1_im) : $signed(matrix_L_inv_1_im); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_57 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_1_re) : $signed(matrix_L_inv_1_re); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_58 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_2_im) : $signed(matrix_L_inv_2_im); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_59 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_2_re) : $signed(matrix_L_inv_2_re); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_60 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_3_im) : $signed(matrix_L_inv_3_im); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_61 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_3_re) : $signed(matrix_L_inv_3_re); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_62 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_4_im) : $signed(matrix_L_inv_4_im); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_63 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_4_re) : $signed(matrix_L_inv_4_re); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_64 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_5_im) : $signed(matrix_L_inv_5_im); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_65 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_5_re) : $signed(matrix_L_inv_5_re); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_66 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_6_im) : $signed(matrix_L_inv_6_im); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_67 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_6_re) : $signed(matrix_L_inv_6_re); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_68 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_7_im) : $signed(matrix_L_inv_7_im); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_69 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_7_re) : $signed(matrix_L_inv_7_re); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_70 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_8_im) : $signed(matrix_L_inv_8_im); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_71 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_8_re) : $signed(matrix_L_inv_8_re); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_72 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_9_im) : $signed(matrix_L_inv_9_im); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [63:0] _GEN_73 = lower_triangular_matrix_inversion_complex_v1_io_valid ? $signed(
    lower_triangular_matrix_inversion_complex_v1_io_matrixOut_9_re) : $signed(matrix_L_inv_9_re); // @[Stap_Main.scala 174:67 175:22 63:39]
  wire [7:0] _GEN_74 = lower_triangular_matrix_inversion_complex_v1_io_valid ? _status_T_1 : status; // @[Stap_Main.scala 174:67 176:16 66:29]
  wire [63:0] _GEN_75 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_0_im) : $signed(matrix_R_inv_0_im); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_76 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_0_re) : $signed(matrix_R_inv_0_re); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_77 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_1_im) : $signed(matrix_R_inv_1_im); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_78 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_1_re) : $signed(matrix_R_inv_1_re); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_79 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_2_im) : $signed(matrix_R_inv_2_im); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_80 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_2_re) : $signed(matrix_R_inv_2_re); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_81 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_3_im) : $signed(matrix_R_inv_3_im); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_82 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_3_re) : $signed(matrix_R_inv_3_re); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_83 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_4_im) : $signed(matrix_R_inv_4_im); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_84 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_4_re) : $signed(matrix_R_inv_4_re); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_85 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_5_im) : $signed(matrix_R_inv_5_im); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_86 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_5_re) : $signed(matrix_R_inv_5_re); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_87 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_6_im) : $signed(matrix_R_inv_6_im); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_88 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_6_re) : $signed(matrix_R_inv_6_re); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_89 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_7_im) : $signed(matrix_R_inv_7_im); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_90 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_7_re) : $signed(matrix_R_inv_7_re); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_91 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_8_im) : $signed(matrix_R_inv_8_im); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_92 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_8_re) : $signed(matrix_R_inv_8_re); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_93 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_9_im) : $signed(matrix_R_inv_9_im); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_94 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_9_re) : $signed(matrix_R_inv_9_re); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_95 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_10_im) : $signed(matrix_R_inv_10_im); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_96 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_10_re) : $signed(matrix_R_inv_10_re); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_97 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_11_im) : $signed(matrix_R_inv_11_im); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_98 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_11_re) : $signed(matrix_R_inv_11_re); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_99 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_12_im) : $signed(matrix_R_inv_12_im); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_100 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_12_re) : $signed(matrix_R_inv_12_re); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_101 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_13_im) : $signed(matrix_R_inv_13_im); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_102 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_13_re) : $signed(matrix_R_inv_13_re); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_103 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_14_im) : $signed(matrix_R_inv_14_im); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_104 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_14_re) : $signed(matrix_R_inv_14_re); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_105 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_15_im) : $signed(matrix_R_inv_15_im); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [63:0] _GEN_106 = matrix_mul_v1_io_valid ? $signed(matrix_mul_v1_io_matrixC_15_re) : $signed(matrix_R_inv_15_re); // @[Stap_Main.scala 201:36 202:22 64:39]
  wire [7:0] _GEN_107 = matrix_mul_v1_io_valid ? _status_T_1 : status; // @[Stap_Main.scala 201:36 203:16 66:29]
  wire [63:0] _GEN_108 = optimal_weight_vector_io_valid ? $signed(optimal_weight_vector_io_matrixOut_0_im) : $signed(
    matrix_w_0_im); // @[Stap_Main.scala 214:44 215:18 65:35]
  wire [63:0] _GEN_109 = optimal_weight_vector_io_valid ? $signed(optimal_weight_vector_io_matrixOut_0_re) : $signed(
    matrix_w_0_re); // @[Stap_Main.scala 214:44 215:18 65:35]
  wire [63:0] _GEN_110 = optimal_weight_vector_io_valid ? $signed(optimal_weight_vector_io_matrixOut_1_im) : $signed(
    matrix_w_1_im); // @[Stap_Main.scala 214:44 215:18 65:35]
  wire [63:0] _GEN_111 = optimal_weight_vector_io_valid ? $signed(optimal_weight_vector_io_matrixOut_1_re) : $signed(
    matrix_w_1_re); // @[Stap_Main.scala 214:44 215:18 65:35]
  wire [63:0] _GEN_112 = optimal_weight_vector_io_valid ? $signed(optimal_weight_vector_io_matrixOut_2_im) : $signed(
    matrix_w_2_im); // @[Stap_Main.scala 214:44 215:18 65:35]
  wire [63:0] _GEN_113 = optimal_weight_vector_io_valid ? $signed(optimal_weight_vector_io_matrixOut_2_re) : $signed(
    matrix_w_2_re); // @[Stap_Main.scala 214:44 215:18 65:35]
  wire [63:0] _GEN_114 = optimal_weight_vector_io_valid ? $signed(optimal_weight_vector_io_matrixOut_3_im) : $signed(
    matrix_w_3_im); // @[Stap_Main.scala 214:44 215:18 65:35]
  wire [63:0] _GEN_115 = optimal_weight_vector_io_valid ? $signed(optimal_weight_vector_io_matrixOut_3_re) : $signed(
    matrix_w_3_re); // @[Stap_Main.scala 214:44 215:18 65:35]
  wire [7:0] _GEN_116 = optimal_weight_vector_io_valid ? _status_T_1 : status; // @[Stap_Main.scala 214:44 216:16 66:29]
  wire [63:0] _GEN_118 = status == 8'ha ? $signed(_GEN_108) : $signed(matrix_w_0_im); // @[Stap_Main.scala 211:33 65:35]
  wire [63:0] _GEN_119 = status == 8'ha ? $signed(_GEN_109) : $signed(matrix_w_0_re); // @[Stap_Main.scala 211:33 65:35]
  wire [63:0] _GEN_120 = status == 8'ha ? $signed(_GEN_110) : $signed(matrix_w_1_im); // @[Stap_Main.scala 211:33 65:35]
  wire [63:0] _GEN_121 = status == 8'ha ? $signed(_GEN_111) : $signed(matrix_w_1_re); // @[Stap_Main.scala 211:33 65:35]
  wire [63:0] _GEN_122 = status == 8'ha ? $signed(_GEN_112) : $signed(matrix_w_2_im); // @[Stap_Main.scala 211:33 65:35]
  wire [63:0] _GEN_123 = status == 8'ha ? $signed(_GEN_113) : $signed(matrix_w_2_re); // @[Stap_Main.scala 211:33 65:35]
  wire [63:0] _GEN_124 = status == 8'ha ? $signed(_GEN_114) : $signed(matrix_w_3_im); // @[Stap_Main.scala 211:33 65:35]
  wire [63:0] _GEN_125 = status == 8'ha ? $signed(_GEN_115) : $signed(matrix_w_3_re); // @[Stap_Main.scala 211:33 65:35]
  wire [7:0] _GEN_126 = status == 8'ha ? _GEN_116 : status; // @[Stap_Main.scala 211:33 66:29]
  wire [7:0] _GEN_168 = status == 8'h9 ? _status_T_1 : _GEN_126; // @[Stap_Main.scala 205:32 210:14]
  wire [63:0] _GEN_169 = status == 8'h9 ? $signed(matrix_w_0_im) : $signed(_GEN_118); // @[Stap_Main.scala 205:32 65:35]
  wire [63:0] _GEN_170 = status == 8'h9 ? $signed(matrix_w_0_re) : $signed(_GEN_119); // @[Stap_Main.scala 205:32 65:35]
  wire [63:0] _GEN_171 = status == 8'h9 ? $signed(matrix_w_1_im) : $signed(_GEN_120); // @[Stap_Main.scala 205:32 65:35]
  wire [63:0] _GEN_172 = status == 8'h9 ? $signed(matrix_w_1_re) : $signed(_GEN_121); // @[Stap_Main.scala 205:32 65:35]
  wire [63:0] _GEN_173 = status == 8'h9 ? $signed(matrix_w_2_im) : $signed(_GEN_122); // @[Stap_Main.scala 205:32 65:35]
  wire [63:0] _GEN_174 = status == 8'h9 ? $signed(matrix_w_2_re) : $signed(_GEN_123); // @[Stap_Main.scala 205:32 65:35]
  wire [63:0] _GEN_175 = status == 8'h9 ? $signed(matrix_w_3_im) : $signed(_GEN_124); // @[Stap_Main.scala 205:32 65:35]
  wire [63:0] _GEN_176 = status == 8'h9 ? $signed(matrix_w_3_re) : $signed(_GEN_125); // @[Stap_Main.scala 205:32 65:35]
  wire [63:0] _GEN_178 = status == 8'h8 ? $signed(_GEN_75) : $signed(matrix_R_inv_0_im); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_179 = status == 8'h8 ? $signed(_GEN_76) : $signed(matrix_R_inv_0_re); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_180 = status == 8'h8 ? $signed(_GEN_77) : $signed(matrix_R_inv_1_im); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_181 = status == 8'h8 ? $signed(_GEN_78) : $signed(matrix_R_inv_1_re); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_182 = status == 8'h8 ? $signed(_GEN_79) : $signed(matrix_R_inv_2_im); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_183 = status == 8'h8 ? $signed(_GEN_80) : $signed(matrix_R_inv_2_re); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_184 = status == 8'h8 ? $signed(_GEN_81) : $signed(matrix_R_inv_3_im); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_185 = status == 8'h8 ? $signed(_GEN_82) : $signed(matrix_R_inv_3_re); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_186 = status == 8'h8 ? $signed(_GEN_83) : $signed(matrix_R_inv_4_im); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_187 = status == 8'h8 ? $signed(_GEN_84) : $signed(matrix_R_inv_4_re); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_188 = status == 8'h8 ? $signed(_GEN_85) : $signed(matrix_R_inv_5_im); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_189 = status == 8'h8 ? $signed(_GEN_86) : $signed(matrix_R_inv_5_re); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_190 = status == 8'h8 ? $signed(_GEN_87) : $signed(matrix_R_inv_6_im); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_191 = status == 8'h8 ? $signed(_GEN_88) : $signed(matrix_R_inv_6_re); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_192 = status == 8'h8 ? $signed(_GEN_89) : $signed(matrix_R_inv_7_im); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_193 = status == 8'h8 ? $signed(_GEN_90) : $signed(matrix_R_inv_7_re); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_194 = status == 8'h8 ? $signed(_GEN_91) : $signed(matrix_R_inv_8_im); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_195 = status == 8'h8 ? $signed(_GEN_92) : $signed(matrix_R_inv_8_re); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_196 = status == 8'h8 ? $signed(_GEN_93) : $signed(matrix_R_inv_9_im); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_197 = status == 8'h8 ? $signed(_GEN_94) : $signed(matrix_R_inv_9_re); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_198 = status == 8'h8 ? $signed(_GEN_95) : $signed(matrix_R_inv_10_im); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_199 = status == 8'h8 ? $signed(_GEN_96) : $signed(matrix_R_inv_10_re); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_200 = status == 8'h8 ? $signed(_GEN_97) : $signed(matrix_R_inv_11_im); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_201 = status == 8'h8 ? $signed(_GEN_98) : $signed(matrix_R_inv_11_re); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_202 = status == 8'h8 ? $signed(_GEN_99) : $signed(matrix_R_inv_12_im); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_203 = status == 8'h8 ? $signed(_GEN_100) : $signed(matrix_R_inv_12_re); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_204 = status == 8'h8 ? $signed(_GEN_101) : $signed(matrix_R_inv_13_im); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_205 = status == 8'h8 ? $signed(_GEN_102) : $signed(matrix_R_inv_13_re); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_206 = status == 8'h8 ? $signed(_GEN_103) : $signed(matrix_R_inv_14_im); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_207 = status == 8'h8 ? $signed(_GEN_104) : $signed(matrix_R_inv_14_re); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_208 = status == 8'h8 ? $signed(_GEN_105) : $signed(matrix_R_inv_15_im); // @[Stap_Main.scala 198:32 64:39]
  wire [63:0] _GEN_209 = status == 8'h8 ? $signed(_GEN_106) : $signed(matrix_R_inv_15_re); // @[Stap_Main.scala 198:32 64:39]
  wire [7:0] _GEN_210 = status == 8'h8 ? _GEN_107 : _GEN_168; // @[Stap_Main.scala 198:32]
  wire [63:0] _GEN_252 = status == 8'h8 ? $signed(matrix_w_0_im) : $signed(_GEN_169); // @[Stap_Main.scala 198:32 65:35]
  wire [63:0] _GEN_253 = status == 8'h8 ? $signed(matrix_w_0_re) : $signed(_GEN_170); // @[Stap_Main.scala 198:32 65:35]
  wire [63:0] _GEN_254 = status == 8'h8 ? $signed(matrix_w_1_im) : $signed(_GEN_171); // @[Stap_Main.scala 198:32 65:35]
  wire [63:0] _GEN_255 = status == 8'h8 ? $signed(matrix_w_1_re) : $signed(_GEN_172); // @[Stap_Main.scala 198:32 65:35]
  wire [63:0] _GEN_256 = status == 8'h8 ? $signed(matrix_w_2_im) : $signed(_GEN_173); // @[Stap_Main.scala 198:32 65:35]
  wire [63:0] _GEN_257 = status == 8'h8 ? $signed(matrix_w_2_re) : $signed(_GEN_174); // @[Stap_Main.scala 198:32 65:35]
  wire [63:0] _GEN_258 = status == 8'h8 ? $signed(matrix_w_3_im) : $signed(_GEN_175); // @[Stap_Main.scala 198:32 65:35]
  wire [63:0] _GEN_259 = status == 8'h8 ? $signed(matrix_w_3_re) : $signed(_GEN_176); // @[Stap_Main.scala 198:32 65:35]
  wire [7:0] _GEN_325 = status == 8'h7 ? _status_T_1 : _GEN_210; // @[Stap_Main.scala 178:32 197:14]
  wire [63:0] _GEN_326 = status == 8'h7 ? $signed(matrix_R_inv_0_im) : $signed(_GEN_178); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_327 = status == 8'h7 ? $signed(matrix_R_inv_0_re) : $signed(_GEN_179); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_328 = status == 8'h7 ? $signed(matrix_R_inv_1_im) : $signed(_GEN_180); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_329 = status == 8'h7 ? $signed(matrix_R_inv_1_re) : $signed(_GEN_181); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_330 = status == 8'h7 ? $signed(matrix_R_inv_2_im) : $signed(_GEN_182); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_331 = status == 8'h7 ? $signed(matrix_R_inv_2_re) : $signed(_GEN_183); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_332 = status == 8'h7 ? $signed(matrix_R_inv_3_im) : $signed(_GEN_184); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_333 = status == 8'h7 ? $signed(matrix_R_inv_3_re) : $signed(_GEN_185); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_334 = status == 8'h7 ? $signed(matrix_R_inv_4_im) : $signed(_GEN_186); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_335 = status == 8'h7 ? $signed(matrix_R_inv_4_re) : $signed(_GEN_187); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_336 = status == 8'h7 ? $signed(matrix_R_inv_5_im) : $signed(_GEN_188); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_337 = status == 8'h7 ? $signed(matrix_R_inv_5_re) : $signed(_GEN_189); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_338 = status == 8'h7 ? $signed(matrix_R_inv_6_im) : $signed(_GEN_190); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_339 = status == 8'h7 ? $signed(matrix_R_inv_6_re) : $signed(_GEN_191); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_340 = status == 8'h7 ? $signed(matrix_R_inv_7_im) : $signed(_GEN_192); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_341 = status == 8'h7 ? $signed(matrix_R_inv_7_re) : $signed(_GEN_193); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_342 = status == 8'h7 ? $signed(matrix_R_inv_8_im) : $signed(_GEN_194); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_343 = status == 8'h7 ? $signed(matrix_R_inv_8_re) : $signed(_GEN_195); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_344 = status == 8'h7 ? $signed(matrix_R_inv_9_im) : $signed(_GEN_196); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_345 = status == 8'h7 ? $signed(matrix_R_inv_9_re) : $signed(_GEN_197); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_346 = status == 8'h7 ? $signed(matrix_R_inv_10_im) : $signed(_GEN_198); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_347 = status == 8'h7 ? $signed(matrix_R_inv_10_re) : $signed(_GEN_199); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_348 = status == 8'h7 ? $signed(matrix_R_inv_11_im) : $signed(_GEN_200); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_349 = status == 8'h7 ? $signed(matrix_R_inv_11_re) : $signed(_GEN_201); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_350 = status == 8'h7 ? $signed(matrix_R_inv_12_im) : $signed(_GEN_202); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_351 = status == 8'h7 ? $signed(matrix_R_inv_12_re) : $signed(_GEN_203); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_352 = status == 8'h7 ? $signed(matrix_R_inv_13_im) : $signed(_GEN_204); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_353 = status == 8'h7 ? $signed(matrix_R_inv_13_re) : $signed(_GEN_205); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_354 = status == 8'h7 ? $signed(matrix_R_inv_14_im) : $signed(_GEN_206); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_355 = status == 8'h7 ? $signed(matrix_R_inv_14_re) : $signed(_GEN_207); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_356 = status == 8'h7 ? $signed(matrix_R_inv_15_im) : $signed(_GEN_208); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_357 = status == 8'h7 ? $signed(matrix_R_inv_15_re) : $signed(_GEN_209); // @[Stap_Main.scala 178:32 64:39]
  wire [63:0] _GEN_399 = status == 8'h7 ? $signed(matrix_w_0_im) : $signed(_GEN_252); // @[Stap_Main.scala 178:32 65:35]
  wire [63:0] _GEN_400 = status == 8'h7 ? $signed(matrix_w_0_re) : $signed(_GEN_253); // @[Stap_Main.scala 178:32 65:35]
  wire [63:0] _GEN_401 = status == 8'h7 ? $signed(matrix_w_1_im) : $signed(_GEN_254); // @[Stap_Main.scala 178:32 65:35]
  wire [63:0] _GEN_402 = status == 8'h7 ? $signed(matrix_w_1_re) : $signed(_GEN_255); // @[Stap_Main.scala 178:32 65:35]
  wire [63:0] _GEN_403 = status == 8'h7 ? $signed(matrix_w_2_im) : $signed(_GEN_256); // @[Stap_Main.scala 178:32 65:35]
  wire [63:0] _GEN_404 = status == 8'h7 ? $signed(matrix_w_2_re) : $signed(_GEN_257); // @[Stap_Main.scala 178:32 65:35]
  wire [63:0] _GEN_405 = status == 8'h7 ? $signed(matrix_w_3_im) : $signed(_GEN_258); // @[Stap_Main.scala 178:32 65:35]
  wire [63:0] _GEN_406 = status == 8'h7 ? $signed(matrix_w_3_re) : $signed(_GEN_259); // @[Stap_Main.scala 178:32 65:35]
  wire [63:0] _GEN_408 = status == 8'h6 ? $signed(_GEN_54) : $signed(matrix_L_inv_0_im); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_409 = status == 8'h6 ? $signed(_GEN_55) : $signed(matrix_L_inv_0_re); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_410 = status == 8'h6 ? $signed(_GEN_56) : $signed(matrix_L_inv_1_im); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_411 = status == 8'h6 ? $signed(_GEN_57) : $signed(matrix_L_inv_1_re); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_412 = status == 8'h6 ? $signed(_GEN_58) : $signed(matrix_L_inv_2_im); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_413 = status == 8'h6 ? $signed(_GEN_59) : $signed(matrix_L_inv_2_re); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_414 = status == 8'h6 ? $signed(_GEN_60) : $signed(matrix_L_inv_3_im); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_415 = status == 8'h6 ? $signed(_GEN_61) : $signed(matrix_L_inv_3_re); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_416 = status == 8'h6 ? $signed(_GEN_62) : $signed(matrix_L_inv_4_im); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_417 = status == 8'h6 ? $signed(_GEN_63) : $signed(matrix_L_inv_4_re); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_418 = status == 8'h6 ? $signed(_GEN_64) : $signed(matrix_L_inv_5_im); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_419 = status == 8'h6 ? $signed(_GEN_65) : $signed(matrix_L_inv_5_re); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_420 = status == 8'h6 ? $signed(_GEN_66) : $signed(matrix_L_inv_6_im); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_421 = status == 8'h6 ? $signed(_GEN_67) : $signed(matrix_L_inv_6_re); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_422 = status == 8'h6 ? $signed(_GEN_68) : $signed(matrix_L_inv_7_im); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_423 = status == 8'h6 ? $signed(_GEN_69) : $signed(matrix_L_inv_7_re); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_424 = status == 8'h6 ? $signed(_GEN_70) : $signed(matrix_L_inv_8_im); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_425 = status == 8'h6 ? $signed(_GEN_71) : $signed(matrix_L_inv_8_re); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_426 = status == 8'h6 ? $signed(_GEN_72) : $signed(matrix_L_inv_9_im); // @[Stap_Main.scala 171:32 63:39]
  wire [63:0] _GEN_427 = status == 8'h6 ? $signed(_GEN_73) : $signed(matrix_L_inv_9_re); // @[Stap_Main.scala 171:32 63:39]
  wire [7:0] _GEN_428 = status == 8'h6 ? _GEN_74 : _GEN_325; // @[Stap_Main.scala 171:32]
  wire [63:0] _GEN_494 = status == 8'h6 ? $signed(matrix_R_inv_0_im) : $signed(_GEN_326); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_495 = status == 8'h6 ? $signed(matrix_R_inv_0_re) : $signed(_GEN_327); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_496 = status == 8'h6 ? $signed(matrix_R_inv_1_im) : $signed(_GEN_328); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_497 = status == 8'h6 ? $signed(matrix_R_inv_1_re) : $signed(_GEN_329); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_498 = status == 8'h6 ? $signed(matrix_R_inv_2_im) : $signed(_GEN_330); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_499 = status == 8'h6 ? $signed(matrix_R_inv_2_re) : $signed(_GEN_331); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_500 = status == 8'h6 ? $signed(matrix_R_inv_3_im) : $signed(_GEN_332); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_501 = status == 8'h6 ? $signed(matrix_R_inv_3_re) : $signed(_GEN_333); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_502 = status == 8'h6 ? $signed(matrix_R_inv_4_im) : $signed(_GEN_334); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_503 = status == 8'h6 ? $signed(matrix_R_inv_4_re) : $signed(_GEN_335); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_504 = status == 8'h6 ? $signed(matrix_R_inv_5_im) : $signed(_GEN_336); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_505 = status == 8'h6 ? $signed(matrix_R_inv_5_re) : $signed(_GEN_337); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_506 = status == 8'h6 ? $signed(matrix_R_inv_6_im) : $signed(_GEN_338); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_507 = status == 8'h6 ? $signed(matrix_R_inv_6_re) : $signed(_GEN_339); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_508 = status == 8'h6 ? $signed(matrix_R_inv_7_im) : $signed(_GEN_340); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_509 = status == 8'h6 ? $signed(matrix_R_inv_7_re) : $signed(_GEN_341); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_510 = status == 8'h6 ? $signed(matrix_R_inv_8_im) : $signed(_GEN_342); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_511 = status == 8'h6 ? $signed(matrix_R_inv_8_re) : $signed(_GEN_343); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_512 = status == 8'h6 ? $signed(matrix_R_inv_9_im) : $signed(_GEN_344); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_513 = status == 8'h6 ? $signed(matrix_R_inv_9_re) : $signed(_GEN_345); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_514 = status == 8'h6 ? $signed(matrix_R_inv_10_im) : $signed(_GEN_346); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_515 = status == 8'h6 ? $signed(matrix_R_inv_10_re) : $signed(_GEN_347); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_516 = status == 8'h6 ? $signed(matrix_R_inv_11_im) : $signed(_GEN_348); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_517 = status == 8'h6 ? $signed(matrix_R_inv_11_re) : $signed(_GEN_349); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_518 = status == 8'h6 ? $signed(matrix_R_inv_12_im) : $signed(_GEN_350); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_519 = status == 8'h6 ? $signed(matrix_R_inv_12_re) : $signed(_GEN_351); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_520 = status == 8'h6 ? $signed(matrix_R_inv_13_im) : $signed(_GEN_352); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_521 = status == 8'h6 ? $signed(matrix_R_inv_13_re) : $signed(_GEN_353); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_522 = status == 8'h6 ? $signed(matrix_R_inv_14_im) : $signed(_GEN_354); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_523 = status == 8'h6 ? $signed(matrix_R_inv_14_re) : $signed(_GEN_355); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_524 = status == 8'h6 ? $signed(matrix_R_inv_15_im) : $signed(_GEN_356); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_525 = status == 8'h6 ? $signed(matrix_R_inv_15_re) : $signed(_GEN_357); // @[Stap_Main.scala 171:32 64:39]
  wire [63:0] _GEN_567 = status == 8'h6 ? $signed(matrix_w_0_im) : $signed(_GEN_399); // @[Stap_Main.scala 171:32 65:35]
  wire [63:0] _GEN_568 = status == 8'h6 ? $signed(matrix_w_0_re) : $signed(_GEN_400); // @[Stap_Main.scala 171:32 65:35]
  wire [63:0] _GEN_569 = status == 8'h6 ? $signed(matrix_w_1_im) : $signed(_GEN_401); // @[Stap_Main.scala 171:32 65:35]
  wire [63:0] _GEN_570 = status == 8'h6 ? $signed(matrix_w_1_re) : $signed(_GEN_402); // @[Stap_Main.scala 171:32 65:35]
  wire [63:0] _GEN_571 = status == 8'h6 ? $signed(matrix_w_2_im) : $signed(_GEN_403); // @[Stap_Main.scala 171:32 65:35]
  wire [63:0] _GEN_572 = status == 8'h6 ? $signed(matrix_w_2_re) : $signed(_GEN_404); // @[Stap_Main.scala 171:32 65:35]
  wire [63:0] _GEN_573 = status == 8'h6 ? $signed(matrix_w_3_im) : $signed(_GEN_405); // @[Stap_Main.scala 171:32 65:35]
  wire [63:0] _GEN_574 = status == 8'h6 ? $signed(matrix_w_3_re) : $signed(_GEN_406); // @[Stap_Main.scala 171:32 65:35]
  wire [7:0] _GEN_596 = status == 8'h5 ? _status_T_1 : _GEN_428; // @[Stap_Main.scala 166:32 170:14]
  wire [63:0] _GEN_597 = status == 8'h5 ? $signed(matrix_L_inv_0_im) : $signed(_GEN_408); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_598 = status == 8'h5 ? $signed(matrix_L_inv_0_re) : $signed(_GEN_409); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_599 = status == 8'h5 ? $signed(matrix_L_inv_1_im) : $signed(_GEN_410); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_600 = status == 8'h5 ? $signed(matrix_L_inv_1_re) : $signed(_GEN_411); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_601 = status == 8'h5 ? $signed(matrix_L_inv_2_im) : $signed(_GEN_412); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_602 = status == 8'h5 ? $signed(matrix_L_inv_2_re) : $signed(_GEN_413); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_603 = status == 8'h5 ? $signed(matrix_L_inv_3_im) : $signed(_GEN_414); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_604 = status == 8'h5 ? $signed(matrix_L_inv_3_re) : $signed(_GEN_415); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_605 = status == 8'h5 ? $signed(matrix_L_inv_4_im) : $signed(_GEN_416); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_606 = status == 8'h5 ? $signed(matrix_L_inv_4_re) : $signed(_GEN_417); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_607 = status == 8'h5 ? $signed(matrix_L_inv_5_im) : $signed(_GEN_418); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_608 = status == 8'h5 ? $signed(matrix_L_inv_5_re) : $signed(_GEN_419); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_609 = status == 8'h5 ? $signed(matrix_L_inv_6_im) : $signed(_GEN_420); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_610 = status == 8'h5 ? $signed(matrix_L_inv_6_re) : $signed(_GEN_421); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_611 = status == 8'h5 ? $signed(matrix_L_inv_7_im) : $signed(_GEN_422); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_612 = status == 8'h5 ? $signed(matrix_L_inv_7_re) : $signed(_GEN_423); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_613 = status == 8'h5 ? $signed(matrix_L_inv_8_im) : $signed(_GEN_424); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_614 = status == 8'h5 ? $signed(matrix_L_inv_8_re) : $signed(_GEN_425); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_615 = status == 8'h5 ? $signed(matrix_L_inv_9_im) : $signed(_GEN_426); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_616 = status == 8'h5 ? $signed(matrix_L_inv_9_re) : $signed(_GEN_427); // @[Stap_Main.scala 166:32 63:39]
  wire [63:0] _GEN_682 = status == 8'h5 ? $signed(matrix_R_inv_0_im) : $signed(_GEN_494); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_683 = status == 8'h5 ? $signed(matrix_R_inv_0_re) : $signed(_GEN_495); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_684 = status == 8'h5 ? $signed(matrix_R_inv_1_im) : $signed(_GEN_496); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_685 = status == 8'h5 ? $signed(matrix_R_inv_1_re) : $signed(_GEN_497); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_686 = status == 8'h5 ? $signed(matrix_R_inv_2_im) : $signed(_GEN_498); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_687 = status == 8'h5 ? $signed(matrix_R_inv_2_re) : $signed(_GEN_499); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_688 = status == 8'h5 ? $signed(matrix_R_inv_3_im) : $signed(_GEN_500); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_689 = status == 8'h5 ? $signed(matrix_R_inv_3_re) : $signed(_GEN_501); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_690 = status == 8'h5 ? $signed(matrix_R_inv_4_im) : $signed(_GEN_502); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_691 = status == 8'h5 ? $signed(matrix_R_inv_4_re) : $signed(_GEN_503); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_692 = status == 8'h5 ? $signed(matrix_R_inv_5_im) : $signed(_GEN_504); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_693 = status == 8'h5 ? $signed(matrix_R_inv_5_re) : $signed(_GEN_505); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_694 = status == 8'h5 ? $signed(matrix_R_inv_6_im) : $signed(_GEN_506); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_695 = status == 8'h5 ? $signed(matrix_R_inv_6_re) : $signed(_GEN_507); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_696 = status == 8'h5 ? $signed(matrix_R_inv_7_im) : $signed(_GEN_508); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_697 = status == 8'h5 ? $signed(matrix_R_inv_7_re) : $signed(_GEN_509); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_698 = status == 8'h5 ? $signed(matrix_R_inv_8_im) : $signed(_GEN_510); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_699 = status == 8'h5 ? $signed(matrix_R_inv_8_re) : $signed(_GEN_511); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_700 = status == 8'h5 ? $signed(matrix_R_inv_9_im) : $signed(_GEN_512); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_701 = status == 8'h5 ? $signed(matrix_R_inv_9_re) : $signed(_GEN_513); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_702 = status == 8'h5 ? $signed(matrix_R_inv_10_im) : $signed(_GEN_514); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_703 = status == 8'h5 ? $signed(matrix_R_inv_10_re) : $signed(_GEN_515); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_704 = status == 8'h5 ? $signed(matrix_R_inv_11_im) : $signed(_GEN_516); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_705 = status == 8'h5 ? $signed(matrix_R_inv_11_re) : $signed(_GEN_517); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_706 = status == 8'h5 ? $signed(matrix_R_inv_12_im) : $signed(_GEN_518); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_707 = status == 8'h5 ? $signed(matrix_R_inv_12_re) : $signed(_GEN_519); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_708 = status == 8'h5 ? $signed(matrix_R_inv_13_im) : $signed(_GEN_520); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_709 = status == 8'h5 ? $signed(matrix_R_inv_13_re) : $signed(_GEN_521); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_710 = status == 8'h5 ? $signed(matrix_R_inv_14_im) : $signed(_GEN_522); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_711 = status == 8'h5 ? $signed(matrix_R_inv_14_re) : $signed(_GEN_523); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_712 = status == 8'h5 ? $signed(matrix_R_inv_15_im) : $signed(_GEN_524); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_713 = status == 8'h5 ? $signed(matrix_R_inv_15_re) : $signed(_GEN_525); // @[Stap_Main.scala 166:32 64:39]
  wire [63:0] _GEN_755 = status == 8'h5 ? $signed(matrix_w_0_im) : $signed(_GEN_567); // @[Stap_Main.scala 166:32 65:35]
  wire [63:0] _GEN_756 = status == 8'h5 ? $signed(matrix_w_0_re) : $signed(_GEN_568); // @[Stap_Main.scala 166:32 65:35]
  wire [63:0] _GEN_757 = status == 8'h5 ? $signed(matrix_w_1_im) : $signed(_GEN_569); // @[Stap_Main.scala 166:32 65:35]
  wire [63:0] _GEN_758 = status == 8'h5 ? $signed(matrix_w_1_re) : $signed(_GEN_570); // @[Stap_Main.scala 166:32 65:35]
  wire [63:0] _GEN_759 = status == 8'h5 ? $signed(matrix_w_2_im) : $signed(_GEN_571); // @[Stap_Main.scala 166:32 65:35]
  wire [63:0] _GEN_760 = status == 8'h5 ? $signed(matrix_w_2_re) : $signed(_GEN_572); // @[Stap_Main.scala 166:32 65:35]
  wire [63:0] _GEN_761 = status == 8'h5 ? $signed(matrix_w_3_im) : $signed(_GEN_573); // @[Stap_Main.scala 166:32 65:35]
  wire [63:0] _GEN_762 = status == 8'h5 ? $signed(matrix_w_3_re) : $signed(_GEN_574); // @[Stap_Main.scala 166:32 65:35]
  wire [63:0] _GEN_764 = status == 8'h4 ? $signed(_GEN_33) : $signed(matrix_L_0_im); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_765 = status == 8'h4 ? $signed(_GEN_34) : $signed(matrix_L_0_re); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_766 = status == 8'h4 ? $signed(_GEN_35) : $signed(matrix_L_1_im); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_767 = status == 8'h4 ? $signed(_GEN_36) : $signed(matrix_L_1_re); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_768 = status == 8'h4 ? $signed(_GEN_37) : $signed(matrix_L_2_im); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_769 = status == 8'h4 ? $signed(_GEN_38) : $signed(matrix_L_2_re); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_770 = status == 8'h4 ? $signed(_GEN_39) : $signed(matrix_L_3_im); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_771 = status == 8'h4 ? $signed(_GEN_40) : $signed(matrix_L_3_re); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_772 = status == 8'h4 ? $signed(_GEN_41) : $signed(matrix_L_4_im); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_773 = status == 8'h4 ? $signed(_GEN_42) : $signed(matrix_L_4_re); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_774 = status == 8'h4 ? $signed(_GEN_43) : $signed(matrix_L_5_im); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_775 = status == 8'h4 ? $signed(_GEN_44) : $signed(matrix_L_5_re); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_776 = status == 8'h4 ? $signed(_GEN_45) : $signed(matrix_L_6_im); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_777 = status == 8'h4 ? $signed(_GEN_46) : $signed(matrix_L_6_re); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_778 = status == 8'h4 ? $signed(_GEN_47) : $signed(matrix_L_7_im); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_779 = status == 8'h4 ? $signed(_GEN_48) : $signed(matrix_L_7_re); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_780 = status == 8'h4 ? $signed(_GEN_49) : $signed(matrix_L_8_im); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_781 = status == 8'h4 ? $signed(_GEN_50) : $signed(matrix_L_8_re); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_782 = status == 8'h4 ? $signed(_GEN_51) : $signed(matrix_L_9_im); // @[Stap_Main.scala 159:32 62:35]
  wire [63:0] _GEN_783 = status == 8'h4 ? $signed(_GEN_52) : $signed(matrix_L_9_re); // @[Stap_Main.scala 159:32 62:35]
  wire [7:0] _GEN_784 = status == 8'h4 ? _GEN_53 : _GEN_596; // @[Stap_Main.scala 159:32]
  wire [63:0] _GEN_806 = status == 8'h4 ? $signed(matrix_L_inv_0_im) : $signed(_GEN_597); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_807 = status == 8'h4 ? $signed(matrix_L_inv_0_re) : $signed(_GEN_598); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_808 = status == 8'h4 ? $signed(matrix_L_inv_1_im) : $signed(_GEN_599); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_809 = status == 8'h4 ? $signed(matrix_L_inv_1_re) : $signed(_GEN_600); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_810 = status == 8'h4 ? $signed(matrix_L_inv_2_im) : $signed(_GEN_601); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_811 = status == 8'h4 ? $signed(matrix_L_inv_2_re) : $signed(_GEN_602); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_812 = status == 8'h4 ? $signed(matrix_L_inv_3_im) : $signed(_GEN_603); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_813 = status == 8'h4 ? $signed(matrix_L_inv_3_re) : $signed(_GEN_604); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_814 = status == 8'h4 ? $signed(matrix_L_inv_4_im) : $signed(_GEN_605); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_815 = status == 8'h4 ? $signed(matrix_L_inv_4_re) : $signed(_GEN_606); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_816 = status == 8'h4 ? $signed(matrix_L_inv_5_im) : $signed(_GEN_607); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_817 = status == 8'h4 ? $signed(matrix_L_inv_5_re) : $signed(_GEN_608); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_818 = status == 8'h4 ? $signed(matrix_L_inv_6_im) : $signed(_GEN_609); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_819 = status == 8'h4 ? $signed(matrix_L_inv_6_re) : $signed(_GEN_610); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_820 = status == 8'h4 ? $signed(matrix_L_inv_7_im) : $signed(_GEN_611); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_821 = status == 8'h4 ? $signed(matrix_L_inv_7_re) : $signed(_GEN_612); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_822 = status == 8'h4 ? $signed(matrix_L_inv_8_im) : $signed(_GEN_613); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_823 = status == 8'h4 ? $signed(matrix_L_inv_8_re) : $signed(_GEN_614); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_824 = status == 8'h4 ? $signed(matrix_L_inv_9_im) : $signed(_GEN_615); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_825 = status == 8'h4 ? $signed(matrix_L_inv_9_re) : $signed(_GEN_616); // @[Stap_Main.scala 159:32 63:39]
  wire [63:0] _GEN_891 = status == 8'h4 ? $signed(matrix_R_inv_0_im) : $signed(_GEN_682); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_892 = status == 8'h4 ? $signed(matrix_R_inv_0_re) : $signed(_GEN_683); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_893 = status == 8'h4 ? $signed(matrix_R_inv_1_im) : $signed(_GEN_684); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_894 = status == 8'h4 ? $signed(matrix_R_inv_1_re) : $signed(_GEN_685); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_895 = status == 8'h4 ? $signed(matrix_R_inv_2_im) : $signed(_GEN_686); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_896 = status == 8'h4 ? $signed(matrix_R_inv_2_re) : $signed(_GEN_687); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_897 = status == 8'h4 ? $signed(matrix_R_inv_3_im) : $signed(_GEN_688); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_898 = status == 8'h4 ? $signed(matrix_R_inv_3_re) : $signed(_GEN_689); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_899 = status == 8'h4 ? $signed(matrix_R_inv_4_im) : $signed(_GEN_690); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_900 = status == 8'h4 ? $signed(matrix_R_inv_4_re) : $signed(_GEN_691); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_901 = status == 8'h4 ? $signed(matrix_R_inv_5_im) : $signed(_GEN_692); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_902 = status == 8'h4 ? $signed(matrix_R_inv_5_re) : $signed(_GEN_693); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_903 = status == 8'h4 ? $signed(matrix_R_inv_6_im) : $signed(_GEN_694); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_904 = status == 8'h4 ? $signed(matrix_R_inv_6_re) : $signed(_GEN_695); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_905 = status == 8'h4 ? $signed(matrix_R_inv_7_im) : $signed(_GEN_696); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_906 = status == 8'h4 ? $signed(matrix_R_inv_7_re) : $signed(_GEN_697); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_907 = status == 8'h4 ? $signed(matrix_R_inv_8_im) : $signed(_GEN_698); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_908 = status == 8'h4 ? $signed(matrix_R_inv_8_re) : $signed(_GEN_699); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_909 = status == 8'h4 ? $signed(matrix_R_inv_9_im) : $signed(_GEN_700); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_910 = status == 8'h4 ? $signed(matrix_R_inv_9_re) : $signed(_GEN_701); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_911 = status == 8'h4 ? $signed(matrix_R_inv_10_im) : $signed(_GEN_702); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_912 = status == 8'h4 ? $signed(matrix_R_inv_10_re) : $signed(_GEN_703); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_913 = status == 8'h4 ? $signed(matrix_R_inv_11_im) : $signed(_GEN_704); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_914 = status == 8'h4 ? $signed(matrix_R_inv_11_re) : $signed(_GEN_705); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_915 = status == 8'h4 ? $signed(matrix_R_inv_12_im) : $signed(_GEN_706); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_916 = status == 8'h4 ? $signed(matrix_R_inv_12_re) : $signed(_GEN_707); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_917 = status == 8'h4 ? $signed(matrix_R_inv_13_im) : $signed(_GEN_708); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_918 = status == 8'h4 ? $signed(matrix_R_inv_13_re) : $signed(_GEN_709); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_919 = status == 8'h4 ? $signed(matrix_R_inv_14_im) : $signed(_GEN_710); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_920 = status == 8'h4 ? $signed(matrix_R_inv_14_re) : $signed(_GEN_711); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_921 = status == 8'h4 ? $signed(matrix_R_inv_15_im) : $signed(_GEN_712); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_922 = status == 8'h4 ? $signed(matrix_R_inv_15_re) : $signed(_GEN_713); // @[Stap_Main.scala 159:32 64:39]
  wire [63:0] _GEN_964 = status == 8'h4 ? $signed(matrix_w_0_im) : $signed(_GEN_755); // @[Stap_Main.scala 159:32 65:35]
  wire [63:0] _GEN_965 = status == 8'h4 ? $signed(matrix_w_0_re) : $signed(_GEN_756); // @[Stap_Main.scala 159:32 65:35]
  wire [63:0] _GEN_966 = status == 8'h4 ? $signed(matrix_w_1_im) : $signed(_GEN_757); // @[Stap_Main.scala 159:32 65:35]
  wire [63:0] _GEN_967 = status == 8'h4 ? $signed(matrix_w_1_re) : $signed(_GEN_758); // @[Stap_Main.scala 159:32 65:35]
  wire [63:0] _GEN_968 = status == 8'h4 ? $signed(matrix_w_2_im) : $signed(_GEN_759); // @[Stap_Main.scala 159:32 65:35]
  wire [63:0] _GEN_969 = status == 8'h4 ? $signed(matrix_w_2_re) : $signed(_GEN_760); // @[Stap_Main.scala 159:32 65:35]
  wire [63:0] _GEN_970 = status == 8'h4 ? $signed(matrix_w_3_im) : $signed(_GEN_761); // @[Stap_Main.scala 159:32 65:35]
  wire [63:0] _GEN_971 = status == 8'h4 ? $signed(matrix_w_3_re) : $signed(_GEN_762); // @[Stap_Main.scala 159:32 65:35]
  wire [7:0] _GEN_1005 = status == 8'h3 ? _status_T_1 : _GEN_784; // @[Stap_Main.scala 154:32 158:14]
  wire [63:0] _GEN_1006 = status == 8'h3 ? $signed(matrix_L_0_im) : $signed(_GEN_764); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1007 = status == 8'h3 ? $signed(matrix_L_0_re) : $signed(_GEN_765); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1008 = status == 8'h3 ? $signed(matrix_L_1_im) : $signed(_GEN_766); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1009 = status == 8'h3 ? $signed(matrix_L_1_re) : $signed(_GEN_767); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1010 = status == 8'h3 ? $signed(matrix_L_2_im) : $signed(_GEN_768); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1011 = status == 8'h3 ? $signed(matrix_L_2_re) : $signed(_GEN_769); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1012 = status == 8'h3 ? $signed(matrix_L_3_im) : $signed(_GEN_770); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1013 = status == 8'h3 ? $signed(matrix_L_3_re) : $signed(_GEN_771); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1014 = status == 8'h3 ? $signed(matrix_L_4_im) : $signed(_GEN_772); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1015 = status == 8'h3 ? $signed(matrix_L_4_re) : $signed(_GEN_773); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1016 = status == 8'h3 ? $signed(matrix_L_5_im) : $signed(_GEN_774); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1017 = status == 8'h3 ? $signed(matrix_L_5_re) : $signed(_GEN_775); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1018 = status == 8'h3 ? $signed(matrix_L_6_im) : $signed(_GEN_776); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1019 = status == 8'h3 ? $signed(matrix_L_6_re) : $signed(_GEN_777); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1020 = status == 8'h3 ? $signed(matrix_L_7_im) : $signed(_GEN_778); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1021 = status == 8'h3 ? $signed(matrix_L_7_re) : $signed(_GEN_779); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1022 = status == 8'h3 ? $signed(matrix_L_8_im) : $signed(_GEN_780); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1023 = status == 8'h3 ? $signed(matrix_L_8_re) : $signed(_GEN_781); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1024 = status == 8'h3 ? $signed(matrix_L_9_im) : $signed(_GEN_782); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1025 = status == 8'h3 ? $signed(matrix_L_9_re) : $signed(_GEN_783); // @[Stap_Main.scala 154:32 62:35]
  wire [63:0] _GEN_1047 = status == 8'h3 ? $signed(matrix_L_inv_0_im) : $signed(_GEN_806); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1048 = status == 8'h3 ? $signed(matrix_L_inv_0_re) : $signed(_GEN_807); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1049 = status == 8'h3 ? $signed(matrix_L_inv_1_im) : $signed(_GEN_808); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1050 = status == 8'h3 ? $signed(matrix_L_inv_1_re) : $signed(_GEN_809); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1051 = status == 8'h3 ? $signed(matrix_L_inv_2_im) : $signed(_GEN_810); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1052 = status == 8'h3 ? $signed(matrix_L_inv_2_re) : $signed(_GEN_811); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1053 = status == 8'h3 ? $signed(matrix_L_inv_3_im) : $signed(_GEN_812); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1054 = status == 8'h3 ? $signed(matrix_L_inv_3_re) : $signed(_GEN_813); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1055 = status == 8'h3 ? $signed(matrix_L_inv_4_im) : $signed(_GEN_814); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1056 = status == 8'h3 ? $signed(matrix_L_inv_4_re) : $signed(_GEN_815); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1057 = status == 8'h3 ? $signed(matrix_L_inv_5_im) : $signed(_GEN_816); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1058 = status == 8'h3 ? $signed(matrix_L_inv_5_re) : $signed(_GEN_817); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1059 = status == 8'h3 ? $signed(matrix_L_inv_6_im) : $signed(_GEN_818); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1060 = status == 8'h3 ? $signed(matrix_L_inv_6_re) : $signed(_GEN_819); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1061 = status == 8'h3 ? $signed(matrix_L_inv_7_im) : $signed(_GEN_820); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1062 = status == 8'h3 ? $signed(matrix_L_inv_7_re) : $signed(_GEN_821); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1063 = status == 8'h3 ? $signed(matrix_L_inv_8_im) : $signed(_GEN_822); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1064 = status == 8'h3 ? $signed(matrix_L_inv_8_re) : $signed(_GEN_823); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1065 = status == 8'h3 ? $signed(matrix_L_inv_9_im) : $signed(_GEN_824); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1066 = status == 8'h3 ? $signed(matrix_L_inv_9_re) : $signed(_GEN_825); // @[Stap_Main.scala 154:32 63:39]
  wire [63:0] _GEN_1132 = status == 8'h3 ? $signed(matrix_R_inv_0_im) : $signed(_GEN_891); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1133 = status == 8'h3 ? $signed(matrix_R_inv_0_re) : $signed(_GEN_892); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1134 = status == 8'h3 ? $signed(matrix_R_inv_1_im) : $signed(_GEN_893); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1135 = status == 8'h3 ? $signed(matrix_R_inv_1_re) : $signed(_GEN_894); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1136 = status == 8'h3 ? $signed(matrix_R_inv_2_im) : $signed(_GEN_895); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1137 = status == 8'h3 ? $signed(matrix_R_inv_2_re) : $signed(_GEN_896); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1138 = status == 8'h3 ? $signed(matrix_R_inv_3_im) : $signed(_GEN_897); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1139 = status == 8'h3 ? $signed(matrix_R_inv_3_re) : $signed(_GEN_898); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1140 = status == 8'h3 ? $signed(matrix_R_inv_4_im) : $signed(_GEN_899); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1141 = status == 8'h3 ? $signed(matrix_R_inv_4_re) : $signed(_GEN_900); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1142 = status == 8'h3 ? $signed(matrix_R_inv_5_im) : $signed(_GEN_901); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1143 = status == 8'h3 ? $signed(matrix_R_inv_5_re) : $signed(_GEN_902); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1144 = status == 8'h3 ? $signed(matrix_R_inv_6_im) : $signed(_GEN_903); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1145 = status == 8'h3 ? $signed(matrix_R_inv_6_re) : $signed(_GEN_904); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1146 = status == 8'h3 ? $signed(matrix_R_inv_7_im) : $signed(_GEN_905); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1147 = status == 8'h3 ? $signed(matrix_R_inv_7_re) : $signed(_GEN_906); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1148 = status == 8'h3 ? $signed(matrix_R_inv_8_im) : $signed(_GEN_907); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1149 = status == 8'h3 ? $signed(matrix_R_inv_8_re) : $signed(_GEN_908); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1150 = status == 8'h3 ? $signed(matrix_R_inv_9_im) : $signed(_GEN_909); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1151 = status == 8'h3 ? $signed(matrix_R_inv_9_re) : $signed(_GEN_910); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1152 = status == 8'h3 ? $signed(matrix_R_inv_10_im) : $signed(_GEN_911); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1153 = status == 8'h3 ? $signed(matrix_R_inv_10_re) : $signed(_GEN_912); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1154 = status == 8'h3 ? $signed(matrix_R_inv_11_im) : $signed(_GEN_913); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1155 = status == 8'h3 ? $signed(matrix_R_inv_11_re) : $signed(_GEN_914); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1156 = status == 8'h3 ? $signed(matrix_R_inv_12_im) : $signed(_GEN_915); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1157 = status == 8'h3 ? $signed(matrix_R_inv_12_re) : $signed(_GEN_916); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1158 = status == 8'h3 ? $signed(matrix_R_inv_13_im) : $signed(_GEN_917); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1159 = status == 8'h3 ? $signed(matrix_R_inv_13_re) : $signed(_GEN_918); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1160 = status == 8'h3 ? $signed(matrix_R_inv_14_im) : $signed(_GEN_919); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1161 = status == 8'h3 ? $signed(matrix_R_inv_14_re) : $signed(_GEN_920); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1162 = status == 8'h3 ? $signed(matrix_R_inv_15_im) : $signed(_GEN_921); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1163 = status == 8'h3 ? $signed(matrix_R_inv_15_re) : $signed(_GEN_922); // @[Stap_Main.scala 154:32 64:39]
  wire [63:0] _GEN_1205 = status == 8'h3 ? $signed(matrix_w_0_im) : $signed(_GEN_964); // @[Stap_Main.scala 154:32 65:35]
  wire [63:0] _GEN_1206 = status == 8'h3 ? $signed(matrix_w_0_re) : $signed(_GEN_965); // @[Stap_Main.scala 154:32 65:35]
  wire [63:0] _GEN_1207 = status == 8'h3 ? $signed(matrix_w_1_im) : $signed(_GEN_966); // @[Stap_Main.scala 154:32 65:35]
  wire [63:0] _GEN_1208 = status == 8'h3 ? $signed(matrix_w_1_re) : $signed(_GEN_967); // @[Stap_Main.scala 154:32 65:35]
  wire [63:0] _GEN_1209 = status == 8'h3 ? $signed(matrix_w_2_im) : $signed(_GEN_968); // @[Stap_Main.scala 154:32 65:35]
  wire [63:0] _GEN_1210 = status == 8'h3 ? $signed(matrix_w_2_re) : $signed(_GEN_969); // @[Stap_Main.scala 154:32 65:35]
  wire [63:0] _GEN_1211 = status == 8'h3 ? $signed(matrix_w_3_im) : $signed(_GEN_970); // @[Stap_Main.scala 154:32 65:35]
  wire [63:0] _GEN_1212 = status == 8'h3 ? $signed(matrix_w_3_re) : $signed(_GEN_971); // @[Stap_Main.scala 154:32 65:35]
  wire [7:0] _GEN_1246 = status == 8'h2 ? _GEN_32 : _GEN_1005; // @[Stap_Main.scala 147:32]
  space_time_steering_vector space_time_steering_vector_unit ( // @[Stap_Main.scala 81:47]
    .clock(space_time_steering_vector_unit_clock),
    .reset(space_time_steering_vector_unit_reset),
    .io_theta(space_time_steering_vector_unit_io_theta),
    .io_psi(space_time_steering_vector_unit_io_psi),
    .io_d(space_time_steering_vector_unit_io_d),
    .io_lambda(space_time_steering_vector_unit_io_lambda),
    .io_v(space_time_steering_vector_unit_io_v),
    .io_T(space_time_steering_vector_unit_io_T),
    .io_matrixOut_0_re(space_time_steering_vector_unit_io_matrixOut_0_re),
    .io_matrixOut_0_im(space_time_steering_vector_unit_io_matrixOut_0_im),
    .io_matrixOut_1_re(space_time_steering_vector_unit_io_matrixOut_1_re),
    .io_matrixOut_1_im(space_time_steering_vector_unit_io_matrixOut_1_im),
    .io_matrixOut_2_re(space_time_steering_vector_unit_io_matrixOut_2_re),
    .io_matrixOut_2_im(space_time_steering_vector_unit_io_matrixOut_2_im),
    .io_matrixOut_3_re(space_time_steering_vector_unit_io_matrixOut_3_re),
    .io_matrixOut_3_im(space_time_steering_vector_unit_io_matrixOut_3_im)
  );
  R_matirx_estimation R_matirx_estimation ( // @[Stap_Main.scala 91:56]
    .clock(R_matirx_estimation_clock),
    .reset(R_matirx_estimation_reset),
    .io_reset(R_matirx_estimation_io_reset),
    .io_ready(R_matirx_estimation_io_ready),
    .io_matrixIn_0_re(R_matirx_estimation_io_matrixIn_0_re),
    .io_matrixIn_0_im(R_matirx_estimation_io_matrixIn_0_im),
    .io_matrixIn_1_re(R_matirx_estimation_io_matrixIn_1_re),
    .io_matrixIn_1_im(R_matirx_estimation_io_matrixIn_1_im),
    .io_matrixIn_2_re(R_matirx_estimation_io_matrixIn_2_re),
    .io_matrixIn_2_im(R_matirx_estimation_io_matrixIn_2_im),
    .io_matrixIn_3_re(R_matirx_estimation_io_matrixIn_3_re),
    .io_matrixIn_3_im(R_matirx_estimation_io_matrixIn_3_im),
    .io_matrixIn_4_re(R_matirx_estimation_io_matrixIn_4_re),
    .io_matrixIn_4_im(R_matirx_estimation_io_matrixIn_4_im),
    .io_matrixIn_5_re(R_matirx_estimation_io_matrixIn_5_re),
    .io_matrixIn_5_im(R_matirx_estimation_io_matrixIn_5_im),
    .io_matrixIn_6_re(R_matirx_estimation_io_matrixIn_6_re),
    .io_matrixIn_6_im(R_matirx_estimation_io_matrixIn_6_im),
    .io_matrixIn_7_re(R_matirx_estimation_io_matrixIn_7_re),
    .io_matrixIn_7_im(R_matirx_estimation_io_matrixIn_7_im),
    .io_matrixOut_0_re(R_matirx_estimation_io_matrixOut_0_re),
    .io_matrixOut_0_im(R_matirx_estimation_io_matrixOut_0_im),
    .io_matrixOut_1_re(R_matirx_estimation_io_matrixOut_1_re),
    .io_matrixOut_1_im(R_matirx_estimation_io_matrixOut_1_im),
    .io_matrixOut_2_re(R_matirx_estimation_io_matrixOut_2_re),
    .io_matrixOut_2_im(R_matirx_estimation_io_matrixOut_2_im),
    .io_matrixOut_3_re(R_matirx_estimation_io_matrixOut_3_re),
    .io_matrixOut_3_im(R_matirx_estimation_io_matrixOut_3_im),
    .io_matrixOut_4_re(R_matirx_estimation_io_matrixOut_4_re),
    .io_matrixOut_4_im(R_matirx_estimation_io_matrixOut_4_im),
    .io_matrixOut_5_re(R_matirx_estimation_io_matrixOut_5_re),
    .io_matrixOut_5_im(R_matirx_estimation_io_matrixOut_5_im),
    .io_matrixOut_6_re(R_matirx_estimation_io_matrixOut_6_re),
    .io_matrixOut_6_im(R_matirx_estimation_io_matrixOut_6_im),
    .io_matrixOut_7_re(R_matirx_estimation_io_matrixOut_7_re),
    .io_matrixOut_7_im(R_matirx_estimation_io_matrixOut_7_im),
    .io_matrixOut_8_re(R_matirx_estimation_io_matrixOut_8_re),
    .io_matrixOut_8_im(R_matirx_estimation_io_matrixOut_8_im),
    .io_matrixOut_9_re(R_matirx_estimation_io_matrixOut_9_re),
    .io_matrixOut_9_im(R_matirx_estimation_io_matrixOut_9_im),
    .io_matrixOut_10_re(R_matirx_estimation_io_matrixOut_10_re),
    .io_matrixOut_10_im(R_matirx_estimation_io_matrixOut_10_im),
    .io_matrixOut_11_re(R_matirx_estimation_io_matrixOut_11_re),
    .io_matrixOut_11_im(R_matirx_estimation_io_matrixOut_11_im),
    .io_matrixOut_12_re(R_matirx_estimation_io_matrixOut_12_re),
    .io_matrixOut_12_im(R_matirx_estimation_io_matrixOut_12_im),
    .io_matrixOut_13_re(R_matirx_estimation_io_matrixOut_13_re),
    .io_matrixOut_13_im(R_matirx_estimation_io_matrixOut_13_im),
    .io_matrixOut_14_re(R_matirx_estimation_io_matrixOut_14_re),
    .io_matrixOut_14_im(R_matirx_estimation_io_matrixOut_14_im),
    .io_matrixOut_15_re(R_matirx_estimation_io_matrixOut_15_re),
    .io_matrixOut_15_im(R_matirx_estimation_io_matrixOut_15_im),
    .io_valid(R_matirx_estimation_io_valid)
  );
  cholesky_v1 cholesky_v1 ( // @[Stap_Main.scala 92:40]
    .clock(cholesky_v1_clock),
    .reset(cholesky_v1_reset),
    .io_reset(cholesky_v1_io_reset),
    .io_ready(cholesky_v1_io_ready),
    .io_matrixIn_0_re(cholesky_v1_io_matrixIn_0_re),
    .io_matrixIn_0_im(cholesky_v1_io_matrixIn_0_im),
    .io_matrixIn_1_re(cholesky_v1_io_matrixIn_1_re),
    .io_matrixIn_1_im(cholesky_v1_io_matrixIn_1_im),
    .io_matrixIn_2_re(cholesky_v1_io_matrixIn_2_re),
    .io_matrixIn_2_im(cholesky_v1_io_matrixIn_2_im),
    .io_matrixIn_3_re(cholesky_v1_io_matrixIn_3_re),
    .io_matrixIn_3_im(cholesky_v1_io_matrixIn_3_im),
    .io_matrixIn_4_re(cholesky_v1_io_matrixIn_4_re),
    .io_matrixIn_4_im(cholesky_v1_io_matrixIn_4_im),
    .io_matrixIn_5_re(cholesky_v1_io_matrixIn_5_re),
    .io_matrixIn_5_im(cholesky_v1_io_matrixIn_5_im),
    .io_matrixIn_6_re(cholesky_v1_io_matrixIn_6_re),
    .io_matrixIn_6_im(cholesky_v1_io_matrixIn_6_im),
    .io_matrixIn_7_re(cholesky_v1_io_matrixIn_7_re),
    .io_matrixIn_7_im(cholesky_v1_io_matrixIn_7_im),
    .io_matrixIn_8_re(cholesky_v1_io_matrixIn_8_re),
    .io_matrixIn_8_im(cholesky_v1_io_matrixIn_8_im),
    .io_matrixIn_9_re(cholesky_v1_io_matrixIn_9_re),
    .io_matrixIn_9_im(cholesky_v1_io_matrixIn_9_im),
    .io_matrixIn_10_re(cholesky_v1_io_matrixIn_10_re),
    .io_matrixIn_10_im(cholesky_v1_io_matrixIn_10_im),
    .io_matrixIn_11_re(cholesky_v1_io_matrixIn_11_re),
    .io_matrixIn_11_im(cholesky_v1_io_matrixIn_11_im),
    .io_matrixIn_12_re(cholesky_v1_io_matrixIn_12_re),
    .io_matrixIn_12_im(cholesky_v1_io_matrixIn_12_im),
    .io_matrixIn_13_re(cholesky_v1_io_matrixIn_13_re),
    .io_matrixIn_13_im(cholesky_v1_io_matrixIn_13_im),
    .io_matrixIn_14_re(cholesky_v1_io_matrixIn_14_re),
    .io_matrixIn_14_im(cholesky_v1_io_matrixIn_14_im),
    .io_matrixIn_15_re(cholesky_v1_io_matrixIn_15_re),
    .io_matrixIn_15_im(cholesky_v1_io_matrixIn_15_im),
    .io_matrixOut_0_re(cholesky_v1_io_matrixOut_0_re),
    .io_matrixOut_0_im(cholesky_v1_io_matrixOut_0_im),
    .io_matrixOut_1_re(cholesky_v1_io_matrixOut_1_re),
    .io_matrixOut_1_im(cholesky_v1_io_matrixOut_1_im),
    .io_matrixOut_2_re(cholesky_v1_io_matrixOut_2_re),
    .io_matrixOut_2_im(cholesky_v1_io_matrixOut_2_im),
    .io_matrixOut_3_re(cholesky_v1_io_matrixOut_3_re),
    .io_matrixOut_3_im(cholesky_v1_io_matrixOut_3_im),
    .io_matrixOut_4_re(cholesky_v1_io_matrixOut_4_re),
    .io_matrixOut_4_im(cholesky_v1_io_matrixOut_4_im),
    .io_matrixOut_5_re(cholesky_v1_io_matrixOut_5_re),
    .io_matrixOut_5_im(cholesky_v1_io_matrixOut_5_im),
    .io_matrixOut_6_re(cholesky_v1_io_matrixOut_6_re),
    .io_matrixOut_6_im(cholesky_v1_io_matrixOut_6_im),
    .io_matrixOut_7_re(cholesky_v1_io_matrixOut_7_re),
    .io_matrixOut_7_im(cholesky_v1_io_matrixOut_7_im),
    .io_matrixOut_8_re(cholesky_v1_io_matrixOut_8_re),
    .io_matrixOut_8_im(cholesky_v1_io_matrixOut_8_im),
    .io_matrixOut_9_re(cholesky_v1_io_matrixOut_9_re),
    .io_matrixOut_9_im(cholesky_v1_io_matrixOut_9_im),
    .io_valid(cholesky_v1_io_valid)
  );
  lower_triangular_matrix_inversion_complex_v1 lower_triangular_matrix_inversion_complex_v1 ( // @[Stap_Main.scala 93:60]
    .clock(lower_triangular_matrix_inversion_complex_v1_clock),
    .reset(lower_triangular_matrix_inversion_complex_v1_reset),
    .io_reset(lower_triangular_matrix_inversion_complex_v1_io_reset),
    .io_ready(lower_triangular_matrix_inversion_complex_v1_io_ready),
    .io_matrixIn_0_re(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_0_re),
    .io_matrixIn_0_im(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_0_im),
    .io_matrixIn_1_re(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_1_re),
    .io_matrixIn_1_im(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_1_im),
    .io_matrixIn_2_re(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_2_re),
    .io_matrixIn_2_im(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_2_im),
    .io_matrixIn_3_re(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_3_re),
    .io_matrixIn_3_im(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_3_im),
    .io_matrixIn_4_re(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_4_re),
    .io_matrixIn_4_im(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_4_im),
    .io_matrixIn_5_re(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_5_re),
    .io_matrixIn_5_im(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_5_im),
    .io_matrixIn_6_re(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_6_re),
    .io_matrixIn_6_im(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_6_im),
    .io_matrixIn_7_re(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_7_re),
    .io_matrixIn_7_im(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_7_im),
    .io_matrixIn_8_re(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_8_re),
    .io_matrixIn_8_im(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_8_im),
    .io_matrixIn_9_re(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_9_re),
    .io_matrixIn_9_im(lower_triangular_matrix_inversion_complex_v1_io_matrixIn_9_im),
    .io_matrixOut_0_re(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_0_re),
    .io_matrixOut_0_im(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_0_im),
    .io_matrixOut_1_re(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_1_re),
    .io_matrixOut_1_im(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_1_im),
    .io_matrixOut_2_re(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_2_re),
    .io_matrixOut_2_im(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_2_im),
    .io_matrixOut_3_re(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_3_re),
    .io_matrixOut_3_im(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_3_im),
    .io_matrixOut_4_re(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_4_re),
    .io_matrixOut_4_im(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_4_im),
    .io_matrixOut_5_re(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_5_re),
    .io_matrixOut_5_im(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_5_im),
    .io_matrixOut_6_re(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_6_re),
    .io_matrixOut_6_im(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_6_im),
    .io_matrixOut_7_re(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_7_re),
    .io_matrixOut_7_im(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_7_im),
    .io_matrixOut_8_re(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_8_re),
    .io_matrixOut_8_im(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_8_im),
    .io_matrixOut_9_re(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_9_re),
    .io_matrixOut_9_im(lower_triangular_matrix_inversion_complex_v1_io_matrixOut_9_im),
    .io_valid(lower_triangular_matrix_inversion_complex_v1_io_valid)
  );
  matrix_mul_v1_2 matrix_mul_v1 ( // @[Stap_Main.scala 94:44]
    .clock(matrix_mul_v1_clock),
    .io_reset(matrix_mul_v1_io_reset),
    .io_ready(matrix_mul_v1_io_ready),
    .io_matrixA_0_re(matrix_mul_v1_io_matrixA_0_re),
    .io_matrixA_0_im(matrix_mul_v1_io_matrixA_0_im),
    .io_matrixA_1_re(matrix_mul_v1_io_matrixA_1_re),
    .io_matrixA_1_im(matrix_mul_v1_io_matrixA_1_im),
    .io_matrixA_2_re(matrix_mul_v1_io_matrixA_2_re),
    .io_matrixA_2_im(matrix_mul_v1_io_matrixA_2_im),
    .io_matrixA_3_re(matrix_mul_v1_io_matrixA_3_re),
    .io_matrixA_3_im(matrix_mul_v1_io_matrixA_3_im),
    .io_matrixA_5_re(matrix_mul_v1_io_matrixA_5_re),
    .io_matrixA_5_im(matrix_mul_v1_io_matrixA_5_im),
    .io_matrixA_6_re(matrix_mul_v1_io_matrixA_6_re),
    .io_matrixA_6_im(matrix_mul_v1_io_matrixA_6_im),
    .io_matrixA_7_re(matrix_mul_v1_io_matrixA_7_re),
    .io_matrixA_7_im(matrix_mul_v1_io_matrixA_7_im),
    .io_matrixA_10_re(matrix_mul_v1_io_matrixA_10_re),
    .io_matrixA_10_im(matrix_mul_v1_io_matrixA_10_im),
    .io_matrixA_11_re(matrix_mul_v1_io_matrixA_11_re),
    .io_matrixA_11_im(matrix_mul_v1_io_matrixA_11_im),
    .io_matrixA_15_re(matrix_mul_v1_io_matrixA_15_re),
    .io_matrixA_15_im(matrix_mul_v1_io_matrixA_15_im),
    .io_matrixB_0_re(matrix_mul_v1_io_matrixB_0_re),
    .io_matrixB_0_im(matrix_mul_v1_io_matrixB_0_im),
    .io_matrixB_4_re(matrix_mul_v1_io_matrixB_4_re),
    .io_matrixB_4_im(matrix_mul_v1_io_matrixB_4_im),
    .io_matrixB_5_re(matrix_mul_v1_io_matrixB_5_re),
    .io_matrixB_5_im(matrix_mul_v1_io_matrixB_5_im),
    .io_matrixB_8_re(matrix_mul_v1_io_matrixB_8_re),
    .io_matrixB_8_im(matrix_mul_v1_io_matrixB_8_im),
    .io_matrixB_9_re(matrix_mul_v1_io_matrixB_9_re),
    .io_matrixB_9_im(matrix_mul_v1_io_matrixB_9_im),
    .io_matrixB_10_re(matrix_mul_v1_io_matrixB_10_re),
    .io_matrixB_10_im(matrix_mul_v1_io_matrixB_10_im),
    .io_matrixB_12_re(matrix_mul_v1_io_matrixB_12_re),
    .io_matrixB_12_im(matrix_mul_v1_io_matrixB_12_im),
    .io_matrixB_13_re(matrix_mul_v1_io_matrixB_13_re),
    .io_matrixB_13_im(matrix_mul_v1_io_matrixB_13_im),
    .io_matrixB_14_re(matrix_mul_v1_io_matrixB_14_re),
    .io_matrixB_14_im(matrix_mul_v1_io_matrixB_14_im),
    .io_matrixB_15_re(matrix_mul_v1_io_matrixB_15_re),
    .io_matrixB_15_im(matrix_mul_v1_io_matrixB_15_im),
    .io_matrixC_0_re(matrix_mul_v1_io_matrixC_0_re),
    .io_matrixC_0_im(matrix_mul_v1_io_matrixC_0_im),
    .io_matrixC_1_re(matrix_mul_v1_io_matrixC_1_re),
    .io_matrixC_1_im(matrix_mul_v1_io_matrixC_1_im),
    .io_matrixC_2_re(matrix_mul_v1_io_matrixC_2_re),
    .io_matrixC_2_im(matrix_mul_v1_io_matrixC_2_im),
    .io_matrixC_3_re(matrix_mul_v1_io_matrixC_3_re),
    .io_matrixC_3_im(matrix_mul_v1_io_matrixC_3_im),
    .io_matrixC_4_re(matrix_mul_v1_io_matrixC_4_re),
    .io_matrixC_4_im(matrix_mul_v1_io_matrixC_4_im),
    .io_matrixC_5_re(matrix_mul_v1_io_matrixC_5_re),
    .io_matrixC_5_im(matrix_mul_v1_io_matrixC_5_im),
    .io_matrixC_6_re(matrix_mul_v1_io_matrixC_6_re),
    .io_matrixC_6_im(matrix_mul_v1_io_matrixC_6_im),
    .io_matrixC_7_re(matrix_mul_v1_io_matrixC_7_re),
    .io_matrixC_7_im(matrix_mul_v1_io_matrixC_7_im),
    .io_matrixC_8_re(matrix_mul_v1_io_matrixC_8_re),
    .io_matrixC_8_im(matrix_mul_v1_io_matrixC_8_im),
    .io_matrixC_9_re(matrix_mul_v1_io_matrixC_9_re),
    .io_matrixC_9_im(matrix_mul_v1_io_matrixC_9_im),
    .io_matrixC_10_re(matrix_mul_v1_io_matrixC_10_re),
    .io_matrixC_10_im(matrix_mul_v1_io_matrixC_10_im),
    .io_matrixC_11_re(matrix_mul_v1_io_matrixC_11_re),
    .io_matrixC_11_im(matrix_mul_v1_io_matrixC_11_im),
    .io_matrixC_12_re(matrix_mul_v1_io_matrixC_12_re),
    .io_matrixC_12_im(matrix_mul_v1_io_matrixC_12_im),
    .io_matrixC_13_re(matrix_mul_v1_io_matrixC_13_re),
    .io_matrixC_13_im(matrix_mul_v1_io_matrixC_13_im),
    .io_matrixC_14_re(matrix_mul_v1_io_matrixC_14_re),
    .io_matrixC_14_im(matrix_mul_v1_io_matrixC_14_im),
    .io_matrixC_15_re(matrix_mul_v1_io_matrixC_15_re),
    .io_matrixC_15_im(matrix_mul_v1_io_matrixC_15_im),
    .io_valid(matrix_mul_v1_io_valid)
  );
  optimal_weight_vector optimal_weight_vector ( // @[Stap_Main.scala 95:60]
    .clock(optimal_weight_vector_clock),
    .reset(optimal_weight_vector_reset),
    .io_reset(optimal_weight_vector_io_reset),
    .io_ready(optimal_weight_vector_io_ready),
    .io_matrixS_0_re(optimal_weight_vector_io_matrixS_0_re),
    .io_matrixS_0_im(optimal_weight_vector_io_matrixS_0_im),
    .io_matrixS_1_re(optimal_weight_vector_io_matrixS_1_re),
    .io_matrixS_1_im(optimal_weight_vector_io_matrixS_1_im),
    .io_matrixS_2_re(optimal_weight_vector_io_matrixS_2_re),
    .io_matrixS_2_im(optimal_weight_vector_io_matrixS_2_im),
    .io_matrixS_3_re(optimal_weight_vector_io_matrixS_3_re),
    .io_matrixS_3_im(optimal_weight_vector_io_matrixS_3_im),
    .io_matrixR_Inv_0_re(optimal_weight_vector_io_matrixR_Inv_0_re),
    .io_matrixR_Inv_0_im(optimal_weight_vector_io_matrixR_Inv_0_im),
    .io_matrixR_Inv_1_re(optimal_weight_vector_io_matrixR_Inv_1_re),
    .io_matrixR_Inv_1_im(optimal_weight_vector_io_matrixR_Inv_1_im),
    .io_matrixR_Inv_2_re(optimal_weight_vector_io_matrixR_Inv_2_re),
    .io_matrixR_Inv_2_im(optimal_weight_vector_io_matrixR_Inv_2_im),
    .io_matrixR_Inv_3_re(optimal_weight_vector_io_matrixR_Inv_3_re),
    .io_matrixR_Inv_3_im(optimal_weight_vector_io_matrixR_Inv_3_im),
    .io_matrixR_Inv_4_re(optimal_weight_vector_io_matrixR_Inv_4_re),
    .io_matrixR_Inv_4_im(optimal_weight_vector_io_matrixR_Inv_4_im),
    .io_matrixR_Inv_5_re(optimal_weight_vector_io_matrixR_Inv_5_re),
    .io_matrixR_Inv_5_im(optimal_weight_vector_io_matrixR_Inv_5_im),
    .io_matrixR_Inv_6_re(optimal_weight_vector_io_matrixR_Inv_6_re),
    .io_matrixR_Inv_6_im(optimal_weight_vector_io_matrixR_Inv_6_im),
    .io_matrixR_Inv_7_re(optimal_weight_vector_io_matrixR_Inv_7_re),
    .io_matrixR_Inv_7_im(optimal_weight_vector_io_matrixR_Inv_7_im),
    .io_matrixR_Inv_8_re(optimal_weight_vector_io_matrixR_Inv_8_re),
    .io_matrixR_Inv_8_im(optimal_weight_vector_io_matrixR_Inv_8_im),
    .io_matrixR_Inv_9_re(optimal_weight_vector_io_matrixR_Inv_9_re),
    .io_matrixR_Inv_9_im(optimal_weight_vector_io_matrixR_Inv_9_im),
    .io_matrixR_Inv_10_re(optimal_weight_vector_io_matrixR_Inv_10_re),
    .io_matrixR_Inv_10_im(optimal_weight_vector_io_matrixR_Inv_10_im),
    .io_matrixR_Inv_11_re(optimal_weight_vector_io_matrixR_Inv_11_re),
    .io_matrixR_Inv_11_im(optimal_weight_vector_io_matrixR_Inv_11_im),
    .io_matrixR_Inv_12_re(optimal_weight_vector_io_matrixR_Inv_12_re),
    .io_matrixR_Inv_12_im(optimal_weight_vector_io_matrixR_Inv_12_im),
    .io_matrixR_Inv_13_re(optimal_weight_vector_io_matrixR_Inv_13_re),
    .io_matrixR_Inv_13_im(optimal_weight_vector_io_matrixR_Inv_13_im),
    .io_matrixR_Inv_14_re(optimal_weight_vector_io_matrixR_Inv_14_re),
    .io_matrixR_Inv_14_im(optimal_weight_vector_io_matrixR_Inv_14_im),
    .io_matrixR_Inv_15_re(optimal_weight_vector_io_matrixR_Inv_15_re),
    .io_matrixR_Inv_15_im(optimal_weight_vector_io_matrixR_Inv_15_im),
    .io_matrixOut_0_re(optimal_weight_vector_io_matrixOut_0_re),
    .io_matrixOut_0_im(optimal_weight_vector_io_matrixOut_0_im),
    .io_matrixOut_1_re(optimal_weight_vector_io_matrixOut_1_re),
    .io_matrixOut_1_im(optimal_weight_vector_io_matrixOut_1_im),
    .io_matrixOut_2_re(optimal_weight_vector_io_matrixOut_2_re),
    .io_matrixOut_2_im(optimal_weight_vector_io_matrixOut_2_im),
    .io_matrixOut_3_re(optimal_weight_vector_io_matrixOut_3_re),
    .io_matrixOut_3_im(optimal_weight_vector_io_matrixOut_3_im),
    .io_valid(optimal_weight_vector_io_valid)
  );
  matirx_conjugate_transpose_1 unit ( // @[Matirx_Conjugate_Transpose.scala 32:22]
    .io_matrixIn_0_re(unit_io_matrixIn_0_re),
    .io_matrixIn_0_im(unit_io_matrixIn_0_im),
    .io_matrixIn_4_re(unit_io_matrixIn_4_re),
    .io_matrixIn_4_im(unit_io_matrixIn_4_im),
    .io_matrixIn_5_re(unit_io_matrixIn_5_re),
    .io_matrixIn_5_im(unit_io_matrixIn_5_im),
    .io_matrixIn_8_re(unit_io_matrixIn_8_re),
    .io_matrixIn_8_im(unit_io_matrixIn_8_im),
    .io_matrixIn_9_re(unit_io_matrixIn_9_re),
    .io_matrixIn_9_im(unit_io_matrixIn_9_im),
    .io_matrixIn_10_re(unit_io_matrixIn_10_re),
    .io_matrixIn_10_im(unit_io_matrixIn_10_im),
    .io_matrixIn_12_re(unit_io_matrixIn_12_re),
    .io_matrixIn_12_im(unit_io_matrixIn_12_im),
    .io_matrixIn_13_re(unit_io_matrixIn_13_re),
    .io_matrixIn_13_im(unit_io_matrixIn_13_im),
    .io_matrixIn_14_re(unit_io_matrixIn_14_re),
    .io_matrixIn_14_im(unit_io_matrixIn_14_im),
    .io_matrixIn_15_re(unit_io_matrixIn_15_re),
    .io_matrixIn_15_im(unit_io_matrixIn_15_im),
    .io_matrixOut_0_re(unit_io_matrixOut_0_re),
    .io_matrixOut_0_im(unit_io_matrixOut_0_im),
    .io_matrixOut_1_re(unit_io_matrixOut_1_re),
    .io_matrixOut_1_im(unit_io_matrixOut_1_im),
    .io_matrixOut_2_re(unit_io_matrixOut_2_re),
    .io_matrixOut_2_im(unit_io_matrixOut_2_im),
    .io_matrixOut_3_re(unit_io_matrixOut_3_re),
    .io_matrixOut_3_im(unit_io_matrixOut_3_im),
    .io_matrixOut_5_re(unit_io_matrixOut_5_re),
    .io_matrixOut_5_im(unit_io_matrixOut_5_im),
    .io_matrixOut_6_re(unit_io_matrixOut_6_re),
    .io_matrixOut_6_im(unit_io_matrixOut_6_im),
    .io_matrixOut_7_re(unit_io_matrixOut_7_re),
    .io_matrixOut_7_im(unit_io_matrixOut_7_im),
    .io_matrixOut_10_re(unit_io_matrixOut_10_re),
    .io_matrixOut_10_im(unit_io_matrixOut_10_im),
    .io_matrixOut_11_re(unit_io_matrixOut_11_re),
    .io_matrixOut_11_im(unit_io_matrixOut_11_im),
    .io_matrixOut_15_re(unit_io_matrixOut_15_re),
    .io_matrixOut_15_im(unit_io_matrixOut_15_im)
  );
  assign io_matrixOut_0_re = matrix_w_0_re; // @[Stap_Main.scala 226:16]
  assign io_matrixOut_0_im = matrix_w_0_im; // @[Stap_Main.scala 226:16]
  assign io_matrixOut_1_re = matrix_w_1_re; // @[Stap_Main.scala 226:16]
  assign io_matrixOut_1_im = matrix_w_1_im; // @[Stap_Main.scala 226:16]
  assign io_matrixOut_2_re = matrix_w_2_re; // @[Stap_Main.scala 226:16]
  assign io_matrixOut_2_im = matrix_w_2_im; // @[Stap_Main.scala 226:16]
  assign io_matrixOut_3_re = matrix_w_3_re; // @[Stap_Main.scala 226:16]
  assign io_matrixOut_3_im = matrix_w_3_im; // @[Stap_Main.scala 226:16]
  assign io_valid = status == 8'hb; // @[Stap_Main.scala 221:15]
  assign io_debug_status = status; // @[Stap_Main.scala 227:19]
  assign io_debug_valid_R_matirx_estimation = R_matirx_estimation_io_valid; // @[Stap_Main.scala 228:38]
  assign io_debug_valid_cholesky_v1 = cholesky_v1_io_valid; // @[Stap_Main.scala 229:30]
  assign io_debug_valid_lower_triangular_matrix_inversion_complex_v1 =
    lower_triangular_matrix_inversion_complex_v1_io_valid; // @[Stap_Main.scala 230:63]
  assign io_debug_valid_matrix_mul_v1 = matrix_mul_v1_io_valid; // @[Stap_Main.scala 231:32]
  assign io_debug_valid_optimal_weight_vector = optimal_weight_vector_io_valid; // @[Stap_Main.scala 232:40]
  assign io_debug_matrix_x_in_0_re = matrix_x_in_0_re; // @[Stap_Main.scala 69:24]
  assign io_debug_matrix_x_in_0_im = matrix_x_in_0_im; // @[Stap_Main.scala 69:24]
  assign io_debug_matrix_x_in_1_re = matrix_x_in_1_re; // @[Stap_Main.scala 69:24]
  assign io_debug_matrix_x_in_1_im = matrix_x_in_1_im; // @[Stap_Main.scala 69:24]
  assign io_debug_matrix_x_in_2_re = matrix_x_in_2_re; // @[Stap_Main.scala 69:24]
  assign io_debug_matrix_x_in_2_im = matrix_x_in_2_im; // @[Stap_Main.scala 69:24]
  assign io_debug_matrix_x_in_3_re = matrix_x_in_3_re; // @[Stap_Main.scala 69:24]
  assign io_debug_matrix_x_in_3_im = matrix_x_in_3_im; // @[Stap_Main.scala 69:24]
  assign io_debug_matrix_x_in_4_re = matrix_x_in_4_re; // @[Stap_Main.scala 69:24]
  assign io_debug_matrix_x_in_4_im = matrix_x_in_4_im; // @[Stap_Main.scala 69:24]
  assign io_debug_matrix_x_in_5_re = matrix_x_in_5_re; // @[Stap_Main.scala 69:24]
  assign io_debug_matrix_x_in_5_im = matrix_x_in_5_im; // @[Stap_Main.scala 69:24]
  assign io_debug_matrix_x_in_6_re = matrix_x_in_6_re; // @[Stap_Main.scala 69:24]
  assign io_debug_matrix_x_in_6_im = matrix_x_in_6_im; // @[Stap_Main.scala 69:24]
  assign io_debug_matrix_x_in_7_re = matrix_x_in_7_re; // @[Stap_Main.scala 69:24]
  assign io_debug_matrix_x_in_7_im = matrix_x_in_7_im; // @[Stap_Main.scala 69:24]
  assign io_debug_matrix_S_0_re = matrix_S_0_re; // @[Stap_Main.scala 70:21]
  assign io_debug_matrix_S_0_im = matrix_S_0_im; // @[Stap_Main.scala 70:21]
  assign io_debug_matrix_S_1_re = matrix_S_1_re; // @[Stap_Main.scala 70:21]
  assign io_debug_matrix_S_1_im = matrix_S_1_im; // @[Stap_Main.scala 70:21]
  assign io_debug_matrix_S_2_re = matrix_S_2_re; // @[Stap_Main.scala 70:21]
  assign io_debug_matrix_S_2_im = matrix_S_2_im; // @[Stap_Main.scala 70:21]
  assign io_debug_matrix_S_3_re = matrix_S_3_re; // @[Stap_Main.scala 70:21]
  assign io_debug_matrix_S_3_im = matrix_S_3_im; // @[Stap_Main.scala 70:21]
  assign io_debug_matrix_R_0_re = matrix_R_0_re; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_0_im = matrix_R_0_im; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_1_re = matrix_R_1_re; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_1_im = matrix_R_1_im; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_2_re = matrix_R_2_re; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_2_im = matrix_R_2_im; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_3_re = matrix_R_3_re; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_3_im = matrix_R_3_im; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_4_re = matrix_R_4_re; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_4_im = matrix_R_4_im; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_5_re = matrix_R_5_re; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_5_im = matrix_R_5_im; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_6_re = matrix_R_6_re; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_6_im = matrix_R_6_im; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_7_re = matrix_R_7_re; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_7_im = matrix_R_7_im; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_8_re = matrix_R_8_re; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_8_im = matrix_R_8_im; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_9_re = matrix_R_9_re; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_9_im = matrix_R_9_im; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_10_re = matrix_R_10_re; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_10_im = matrix_R_10_im; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_11_re = matrix_R_11_re; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_11_im = matrix_R_11_im; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_12_re = matrix_R_12_re; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_12_im = matrix_R_12_im; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_13_re = matrix_R_13_re; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_13_im = matrix_R_13_im; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_14_re = matrix_R_14_re; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_14_im = matrix_R_14_im; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_15_re = matrix_R_15_re; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_R_15_im = matrix_R_15_im; // @[Stap_Main.scala 71:21]
  assign io_debug_matrix_L_0_re = matrix_L_0_re; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_0_im = matrix_L_0_im; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_1_re = matrix_L_1_re; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_1_im = matrix_L_1_im; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_2_re = matrix_L_2_re; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_2_im = matrix_L_2_im; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_3_re = matrix_L_3_re; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_3_im = matrix_L_3_im; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_4_re = matrix_L_4_re; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_4_im = matrix_L_4_im; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_5_re = matrix_L_5_re; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_5_im = matrix_L_5_im; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_6_re = matrix_L_6_re; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_6_im = matrix_L_6_im; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_7_re = matrix_L_7_re; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_7_im = matrix_L_7_im; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_8_re = matrix_L_8_re; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_8_im = matrix_L_8_im; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_9_re = matrix_L_9_re; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_9_im = matrix_L_9_im; // @[Stap_Main.scala 72:21]
  assign io_debug_matrix_L_inv_0_re = matrix_L_inv_0_re; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_0_im = matrix_L_inv_0_im; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_1_re = matrix_L_inv_1_re; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_1_im = matrix_L_inv_1_im; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_2_re = matrix_L_inv_2_re; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_2_im = matrix_L_inv_2_im; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_3_re = matrix_L_inv_3_re; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_3_im = matrix_L_inv_3_im; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_4_re = matrix_L_inv_4_re; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_4_im = matrix_L_inv_4_im; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_5_re = matrix_L_inv_5_re; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_5_im = matrix_L_inv_5_im; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_6_re = matrix_L_inv_6_re; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_6_im = matrix_L_inv_6_im; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_7_re = matrix_L_inv_7_re; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_7_im = matrix_L_inv_7_im; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_8_re = matrix_L_inv_8_re; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_8_im = matrix_L_inv_8_im; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_9_re = matrix_L_inv_9_re; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_L_inv_9_im = matrix_L_inv_9_im; // @[Stap_Main.scala 73:25]
  assign io_debug_matrix_R_inv_0_re = matrix_R_inv_0_re; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_0_im = matrix_R_inv_0_im; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_1_re = matrix_R_inv_1_re; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_1_im = matrix_R_inv_1_im; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_2_re = matrix_R_inv_2_re; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_2_im = matrix_R_inv_2_im; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_3_re = matrix_R_inv_3_re; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_3_im = matrix_R_inv_3_im; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_4_re = matrix_R_inv_4_re; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_4_im = matrix_R_inv_4_im; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_5_re = matrix_R_inv_5_re; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_5_im = matrix_R_inv_5_im; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_6_re = matrix_R_inv_6_re; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_6_im = matrix_R_inv_6_im; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_7_re = matrix_R_inv_7_re; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_7_im = matrix_R_inv_7_im; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_8_re = matrix_R_inv_8_re; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_8_im = matrix_R_inv_8_im; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_9_re = matrix_R_inv_9_re; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_9_im = matrix_R_inv_9_im; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_10_re = matrix_R_inv_10_re; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_10_im = matrix_R_inv_10_im; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_11_re = matrix_R_inv_11_re; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_11_im = matrix_R_inv_11_im; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_12_re = matrix_R_inv_12_re; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_12_im = matrix_R_inv_12_im; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_13_re = matrix_R_inv_13_re; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_13_im = matrix_R_inv_13_im; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_14_re = matrix_R_inv_14_re; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_14_im = matrix_R_inv_14_im; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_15_re = matrix_R_inv_15_re; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_R_inv_15_im = matrix_R_inv_15_im; // @[Stap_Main.scala 74:25]
  assign io_debug_matrix_w_0_re = matrix_w_0_re; // @[Stap_Main.scala 75:21]
  assign io_debug_matrix_w_0_im = matrix_w_0_im; // @[Stap_Main.scala 75:21]
  assign io_debug_matrix_w_1_re = matrix_w_1_re; // @[Stap_Main.scala 75:21]
  assign io_debug_matrix_w_1_im = matrix_w_1_im; // @[Stap_Main.scala 75:21]
  assign io_debug_matrix_w_2_re = matrix_w_2_re; // @[Stap_Main.scala 75:21]
  assign io_debug_matrix_w_2_im = matrix_w_2_im; // @[Stap_Main.scala 75:21]
  assign io_debug_matrix_w_3_re = matrix_w_3_re; // @[Stap_Main.scala 75:21]
  assign io_debug_matrix_w_3_im = matrix_w_3_im; // @[Stap_Main.scala 75:21]
  assign space_time_steering_vector_unit_clock = clock;
  assign space_time_steering_vector_unit_reset = reset;
  assign space_time_steering_vector_unit_io_theta = io_theta; // @[Stap_Main.scala 82:44]
  assign space_time_steering_vector_unit_io_psi = io_psi; // @[Stap_Main.scala 83:42]
  assign space_time_steering_vector_unit_io_d = io_d; // @[Stap_Main.scala 84:40]
  assign space_time_steering_vector_unit_io_lambda = io_lambda; // @[Stap_Main.scala 85:45]
  assign space_time_steering_vector_unit_io_v = io_v; // @[Stap_Main.scala 86:40]
  assign space_time_steering_vector_unit_io_T = io_T; // @[Stap_Main.scala 87:40]
  assign R_matirx_estimation_clock = clock;
  assign R_matirx_estimation_reset = reset;
  assign R_matirx_estimation_io_reset = io_reset; // @[Stap_Main.scala 96:32]
  assign R_matirx_estimation_io_ready = status == 8'h1; // @[Stap_Main.scala 142:17]
  assign R_matirx_estimation_io_matrixIn_0_re = matrix_x_in_0_re; // @[Stap_Main.scala 142:26 145:39]
  assign R_matirx_estimation_io_matrixIn_0_im = matrix_x_in_0_im; // @[Stap_Main.scala 142:26 145:39]
  assign R_matirx_estimation_io_matrixIn_1_re = matrix_x_in_1_re; // @[Stap_Main.scala 142:26 145:39]
  assign R_matirx_estimation_io_matrixIn_1_im = matrix_x_in_1_im; // @[Stap_Main.scala 142:26 145:39]
  assign R_matirx_estimation_io_matrixIn_2_re = matrix_x_in_2_re; // @[Stap_Main.scala 142:26 145:39]
  assign R_matirx_estimation_io_matrixIn_2_im = matrix_x_in_2_im; // @[Stap_Main.scala 142:26 145:39]
  assign R_matirx_estimation_io_matrixIn_3_re = matrix_x_in_3_re; // @[Stap_Main.scala 142:26 145:39]
  assign R_matirx_estimation_io_matrixIn_3_im = matrix_x_in_3_im; // @[Stap_Main.scala 142:26 145:39]
  assign R_matirx_estimation_io_matrixIn_4_re = matrix_x_in_4_re; // @[Stap_Main.scala 142:26 145:39]
  assign R_matirx_estimation_io_matrixIn_4_im = matrix_x_in_4_im; // @[Stap_Main.scala 142:26 145:39]
  assign R_matirx_estimation_io_matrixIn_5_re = matrix_x_in_5_re; // @[Stap_Main.scala 142:26 145:39]
  assign R_matirx_estimation_io_matrixIn_5_im = matrix_x_in_5_im; // @[Stap_Main.scala 142:26 145:39]
  assign R_matirx_estimation_io_matrixIn_6_re = matrix_x_in_6_re; // @[Stap_Main.scala 142:26 145:39]
  assign R_matirx_estimation_io_matrixIn_6_im = matrix_x_in_6_im; // @[Stap_Main.scala 142:26 145:39]
  assign R_matirx_estimation_io_matrixIn_7_re = matrix_x_in_7_re; // @[Stap_Main.scala 142:26 145:39]
  assign R_matirx_estimation_io_matrixIn_7_im = matrix_x_in_7_im; // @[Stap_Main.scala 142:26 145:39]
  assign cholesky_v1_clock = clock;
  assign cholesky_v1_reset = reset;
  assign cholesky_v1_io_reset = io_reset; // @[Stap_Main.scala 99:24]
  assign cholesky_v1_io_ready = status == 8'h3; // @[Stap_Main.scala 154:23]
  assign cholesky_v1_io_matrixIn_0_re = matrix_R_0_re; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_0_im = matrix_R_0_im; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_1_re = matrix_R_1_re; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_1_im = matrix_R_1_im; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_2_re = matrix_R_2_re; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_2_im = matrix_R_2_im; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_3_re = matrix_R_3_re; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_3_im = matrix_R_3_im; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_4_re = matrix_R_4_re; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_4_im = matrix_R_4_im; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_5_re = matrix_R_5_re; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_5_im = matrix_R_5_im; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_6_re = matrix_R_6_re; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_6_im = matrix_R_6_im; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_7_re = matrix_R_7_re; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_7_im = matrix_R_7_im; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_8_re = matrix_R_8_re; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_8_im = matrix_R_8_im; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_9_re = matrix_R_9_re; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_9_im = matrix_R_9_im; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_10_re = matrix_R_10_re; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_10_im = matrix_R_10_im; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_11_re = matrix_R_11_re; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_11_im = matrix_R_11_im; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_12_re = matrix_R_12_re; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_12_im = matrix_R_12_im; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_13_re = matrix_R_13_re; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_13_im = matrix_R_13_im; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_14_re = matrix_R_14_re; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_14_im = matrix_R_14_im; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_15_re = matrix_R_15_re; // @[Stap_Main.scala 154:32 157:31]
  assign cholesky_v1_io_matrixIn_15_im = matrix_R_15_im; // @[Stap_Main.scala 154:32 157:31]
  assign lower_triangular_matrix_inversion_complex_v1_clock = clock;
  assign lower_triangular_matrix_inversion_complex_v1_reset = reset;
  assign lower_triangular_matrix_inversion_complex_v1_io_reset = io_reset; // @[Stap_Main.scala 102:57]
  assign lower_triangular_matrix_inversion_complex_v1_io_ready = status == 8'h5; // @[Stap_Main.scala 166:23]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_0_re = matrix_L_0_re; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_0_im = matrix_L_0_im; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_1_re = matrix_L_1_re; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_1_im = matrix_L_1_im; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_2_re = matrix_L_2_re; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_2_im = matrix_L_2_im; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_3_re = matrix_L_3_re; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_3_im = matrix_L_3_im; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_4_re = matrix_L_4_re; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_4_im = matrix_L_4_im; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_5_re = matrix_L_5_re; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_5_im = matrix_L_5_im; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_6_re = matrix_L_6_re; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_6_im = matrix_L_6_im; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_7_re = matrix_L_7_re; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_7_im = matrix_L_7_im; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_8_re = matrix_L_8_re; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_8_im = matrix_L_8_im; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_9_re = matrix_L_9_re; // @[Stap_Main.scala 166:32 169:64]
  assign lower_triangular_matrix_inversion_complex_v1_io_matrixIn_9_im = matrix_L_9_im; // @[Stap_Main.scala 166:32 169:64]
  assign matrix_mul_v1_clock = clock;
  assign matrix_mul_v1_io_reset = io_reset; // @[Stap_Main.scala 105:26]
  assign matrix_mul_v1_io_ready = status == 8'h7; // @[Stap_Main.scala 178:23]
  assign matrix_mul_v1_io_matrixA_0_re = unit_io_matrixOut_0_re; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_0_im = unit_io_matrixOut_0_im; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_1_re = unit_io_matrixOut_1_re; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_1_im = unit_io_matrixOut_1_im; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_2_re = unit_io_matrixOut_2_re; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_2_im = unit_io_matrixOut_2_im; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_3_re = unit_io_matrixOut_3_re; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_3_im = unit_io_matrixOut_3_im; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_5_re = unit_io_matrixOut_5_re; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_5_im = unit_io_matrixOut_5_im; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_6_re = unit_io_matrixOut_6_re; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_6_im = unit_io_matrixOut_6_im; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_7_re = unit_io_matrixOut_7_re; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_7_im = unit_io_matrixOut_7_im; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_10_re = unit_io_matrixOut_10_re; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_10_im = unit_io_matrixOut_10_im; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_11_re = unit_io_matrixOut_11_re; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_11_im = unit_io_matrixOut_11_im; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_15_re = unit_io_matrixOut_15_re; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixA_15_im = unit_io_matrixOut_15_im; // @[Stap_Main.scala 178:32 195:32]
  assign matrix_mul_v1_io_matrixB_0_re = matrix_L_inv_0_re; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_0_im = matrix_L_inv_0_im; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_4_re = matrix_L_inv_1_re; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_4_im = matrix_L_inv_1_im; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_5_re = matrix_L_inv_2_re; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_5_im = matrix_L_inv_2_im; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_8_re = matrix_L_inv_3_re; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_8_im = matrix_L_inv_3_im; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_9_re = matrix_L_inv_4_re; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_9_im = matrix_L_inv_4_im; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_10_re = matrix_L_inv_5_re; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_10_im = matrix_L_inv_5_im; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_12_re = matrix_L_inv_6_re; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_12_im = matrix_L_inv_6_im; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_13_re = matrix_L_inv_7_re; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_13_im = matrix_L_inv_7_im; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_14_re = matrix_L_inv_8_re; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_14_im = matrix_L_inv_8_im; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_15_re = matrix_L_inv_9_re; // @[Stap_Main.scala 180:31 186:38]
  assign matrix_mul_v1_io_matrixB_15_im = matrix_L_inv_9_im; // @[Stap_Main.scala 180:31 186:38]
  assign optimal_weight_vector_clock = clock;
  assign optimal_weight_vector_reset = reset;
  assign optimal_weight_vector_io_reset = io_reset; // @[Stap_Main.scala 109:34]
  assign optimal_weight_vector_io_ready = status == 8'h9; // @[Stap_Main.scala 205:23]
  assign optimal_weight_vector_io_matrixS_0_re = matrix_S_0_re; // @[Stap_Main.scala 205:32 208:40]
  assign optimal_weight_vector_io_matrixS_0_im = matrix_S_0_im; // @[Stap_Main.scala 205:32 208:40]
  assign optimal_weight_vector_io_matrixS_1_re = matrix_S_1_re; // @[Stap_Main.scala 205:32 208:40]
  assign optimal_weight_vector_io_matrixS_1_im = matrix_S_1_im; // @[Stap_Main.scala 205:32 208:40]
  assign optimal_weight_vector_io_matrixS_2_re = matrix_S_2_re; // @[Stap_Main.scala 205:32 208:40]
  assign optimal_weight_vector_io_matrixS_2_im = matrix_S_2_im; // @[Stap_Main.scala 205:32 208:40]
  assign optimal_weight_vector_io_matrixS_3_re = matrix_S_3_re; // @[Stap_Main.scala 205:32 208:40]
  assign optimal_weight_vector_io_matrixS_3_im = matrix_S_3_im; // @[Stap_Main.scala 205:32 208:40]
  assign optimal_weight_vector_io_matrixR_Inv_0_re = matrix_R_inv_0_re; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_0_im = matrix_R_inv_0_im; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_1_re = matrix_R_inv_1_re; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_1_im = matrix_R_inv_1_im; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_2_re = matrix_R_inv_2_re; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_2_im = matrix_R_inv_2_im; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_3_re = matrix_R_inv_3_re; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_3_im = matrix_R_inv_3_im; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_4_re = matrix_R_inv_4_re; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_4_im = matrix_R_inv_4_im; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_5_re = matrix_R_inv_5_re; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_5_im = matrix_R_inv_5_im; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_6_re = matrix_R_inv_6_re; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_6_im = matrix_R_inv_6_im; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_7_re = matrix_R_inv_7_re; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_7_im = matrix_R_inv_7_im; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_8_re = matrix_R_inv_8_re; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_8_im = matrix_R_inv_8_im; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_9_re = matrix_R_inv_9_re; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_9_im = matrix_R_inv_9_im; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_10_re = matrix_R_inv_10_re; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_10_im = matrix_R_inv_10_im; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_11_re = matrix_R_inv_11_re; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_11_im = matrix_R_inv_11_im; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_12_re = matrix_R_inv_12_re; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_12_im = matrix_R_inv_12_im; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_13_re = matrix_R_inv_13_re; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_13_im = matrix_R_inv_13_im; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_14_re = matrix_R_inv_14_re; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_14_im = matrix_R_inv_14_im; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_15_re = matrix_R_inv_15_re; // @[Stap_Main.scala 205:32 209:44]
  assign optimal_weight_vector_io_matrixR_Inv_15_im = matrix_R_inv_15_im; // @[Stap_Main.scala 205:32 209:44]
  assign unit_io_matrixIn_0_re = matrix_L_inv_0_re; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_0_im = matrix_L_inv_0_im; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_4_re = matrix_L_inv_1_re; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_4_im = matrix_L_inv_1_im; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_5_re = matrix_L_inv_2_re; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_5_im = matrix_L_inv_2_im; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_8_re = matrix_L_inv_3_re; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_8_im = matrix_L_inv_3_im; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_9_re = matrix_L_inv_4_re; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_9_im = matrix_L_inv_4_im; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_10_re = matrix_L_inv_5_re; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_10_im = matrix_L_inv_5_im; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_12_re = matrix_L_inv_6_re; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_12_im = matrix_L_inv_6_im; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_13_re = matrix_L_inv_7_re; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_13_im = matrix_L_inv_7_im; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_14_re = matrix_L_inv_8_re; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_14_im = matrix_L_inv_8_im; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_15_re = matrix_L_inv_9_re; // @[Stap_Main.scala 180:31 186:38]
  assign unit_io_matrixIn_15_im = matrix_L_inv_9_im; // @[Stap_Main.scala 180:31 186:38]
  always @(posedge clock) begin
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_x_in_0_re <= 64'sh0; // @[Stap_Main.scala 117:25]
    end else if (io_ready) begin // @[Stap_Main.scala 137:24]
      matrix_x_in_0_re <= io_matrixIn_0_re; // @[Stap_Main.scala 139:17]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_x_in_0_im <= 64'sh0; // @[Stap_Main.scala 118:25]
    end else if (io_ready) begin // @[Stap_Main.scala 137:24]
      matrix_x_in_0_im <= io_matrixIn_0_im; // @[Stap_Main.scala 139:17]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_x_in_1_re <= 64'sh0; // @[Stap_Main.scala 117:25]
    end else if (io_ready) begin // @[Stap_Main.scala 137:24]
      matrix_x_in_1_re <= io_matrixIn_1_re; // @[Stap_Main.scala 139:17]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_x_in_1_im <= 64'sh0; // @[Stap_Main.scala 118:25]
    end else if (io_ready) begin // @[Stap_Main.scala 137:24]
      matrix_x_in_1_im <= io_matrixIn_1_im; // @[Stap_Main.scala 139:17]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_x_in_2_re <= 64'sh0; // @[Stap_Main.scala 117:25]
    end else if (io_ready) begin // @[Stap_Main.scala 137:24]
      matrix_x_in_2_re <= io_matrixIn_2_re; // @[Stap_Main.scala 139:17]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_x_in_2_im <= 64'sh0; // @[Stap_Main.scala 118:25]
    end else if (io_ready) begin // @[Stap_Main.scala 137:24]
      matrix_x_in_2_im <= io_matrixIn_2_im; // @[Stap_Main.scala 139:17]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_x_in_3_re <= 64'sh0; // @[Stap_Main.scala 117:25]
    end else if (io_ready) begin // @[Stap_Main.scala 137:24]
      matrix_x_in_3_re <= io_matrixIn_3_re; // @[Stap_Main.scala 139:17]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_x_in_3_im <= 64'sh0; // @[Stap_Main.scala 118:25]
    end else if (io_ready) begin // @[Stap_Main.scala 137:24]
      matrix_x_in_3_im <= io_matrixIn_3_im; // @[Stap_Main.scala 139:17]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_x_in_4_re <= 64'sh0; // @[Stap_Main.scala 117:25]
    end else if (io_ready) begin // @[Stap_Main.scala 137:24]
      matrix_x_in_4_re <= io_matrixIn_4_re; // @[Stap_Main.scala 139:17]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_x_in_4_im <= 64'sh0; // @[Stap_Main.scala 118:25]
    end else if (io_ready) begin // @[Stap_Main.scala 137:24]
      matrix_x_in_4_im <= io_matrixIn_4_im; // @[Stap_Main.scala 139:17]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_x_in_5_re <= 64'sh0; // @[Stap_Main.scala 117:25]
    end else if (io_ready) begin // @[Stap_Main.scala 137:24]
      matrix_x_in_5_re <= io_matrixIn_5_re; // @[Stap_Main.scala 139:17]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_x_in_5_im <= 64'sh0; // @[Stap_Main.scala 118:25]
    end else if (io_ready) begin // @[Stap_Main.scala 137:24]
      matrix_x_in_5_im <= io_matrixIn_5_im; // @[Stap_Main.scala 139:17]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_x_in_6_re <= 64'sh0; // @[Stap_Main.scala 117:25]
    end else if (io_ready) begin // @[Stap_Main.scala 137:24]
      matrix_x_in_6_re <= io_matrixIn_6_re; // @[Stap_Main.scala 139:17]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_x_in_6_im <= 64'sh0; // @[Stap_Main.scala 118:25]
    end else if (io_ready) begin // @[Stap_Main.scala 137:24]
      matrix_x_in_6_im <= io_matrixIn_6_im; // @[Stap_Main.scala 139:17]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_x_in_7_re <= 64'sh0; // @[Stap_Main.scala 117:25]
    end else if (io_ready) begin // @[Stap_Main.scala 137:24]
      matrix_x_in_7_re <= io_matrixIn_7_re; // @[Stap_Main.scala 139:17]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_x_in_7_im <= 64'sh0; // @[Stap_Main.scala 118:25]
    end else if (io_ready) begin // @[Stap_Main.scala 137:24]
      matrix_x_in_7_im <= io_matrixIn_7_im; // @[Stap_Main.scala 139:17]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_S_0_re <= 64'sh0; // @[Stap_Main.scala 121:22]
    end else begin
      matrix_S_0_re <= space_time_steering_vector_unit_io_matrixOut_0_re; // @[Stap_Main.scala 88:12]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_S_0_im <= 64'sh0; // @[Stap_Main.scala 122:22]
    end else begin
      matrix_S_0_im <= space_time_steering_vector_unit_io_matrixOut_0_im; // @[Stap_Main.scala 88:12]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_S_1_re <= 64'sh0; // @[Stap_Main.scala 121:22]
    end else begin
      matrix_S_1_re <= space_time_steering_vector_unit_io_matrixOut_1_re; // @[Stap_Main.scala 88:12]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_S_1_im <= 64'sh0; // @[Stap_Main.scala 122:22]
    end else begin
      matrix_S_1_im <= space_time_steering_vector_unit_io_matrixOut_1_im; // @[Stap_Main.scala 88:12]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_S_2_re <= 64'sh0; // @[Stap_Main.scala 121:22]
    end else begin
      matrix_S_2_re <= space_time_steering_vector_unit_io_matrixOut_2_re; // @[Stap_Main.scala 88:12]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_S_2_im <= 64'sh0; // @[Stap_Main.scala 122:22]
    end else begin
      matrix_S_2_im <= space_time_steering_vector_unit_io_matrixOut_2_im; // @[Stap_Main.scala 88:12]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_S_3_re <= 64'sh0; // @[Stap_Main.scala 121:22]
    end else begin
      matrix_S_3_re <= space_time_steering_vector_unit_io_matrixOut_3_re; // @[Stap_Main.scala 88:12]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_S_3_im <= 64'sh0; // @[Stap_Main.scala 122:22]
    end else begin
      matrix_S_3_im <= space_time_steering_vector_unit_io_matrixOut_3_im; // @[Stap_Main.scala 88:12]
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_0_re <= 64'sh0; // @[Stap_Main.scala 127:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_0_re <= _GEN_1;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_0_im <= 64'sh0; // @[Stap_Main.scala 128:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_0_im <= _GEN_0;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_1_re <= 64'sh0; // @[Stap_Main.scala 127:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_1_re <= _GEN_3;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_1_im <= 64'sh0; // @[Stap_Main.scala 128:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_1_im <= _GEN_2;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_2_re <= 64'sh0; // @[Stap_Main.scala 127:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_2_re <= _GEN_5;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_2_im <= 64'sh0; // @[Stap_Main.scala 128:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_2_im <= _GEN_4;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_3_re <= 64'sh0; // @[Stap_Main.scala 127:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_3_re <= _GEN_7;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_3_im <= 64'sh0; // @[Stap_Main.scala 128:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_3_im <= _GEN_6;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_4_re <= 64'sh0; // @[Stap_Main.scala 127:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_4_re <= _GEN_9;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_4_im <= 64'sh0; // @[Stap_Main.scala 128:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_4_im <= _GEN_8;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_5_re <= 64'sh0; // @[Stap_Main.scala 127:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_5_re <= _GEN_11;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_5_im <= 64'sh0; // @[Stap_Main.scala 128:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_5_im <= _GEN_10;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_6_re <= 64'sh0; // @[Stap_Main.scala 127:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_6_re <= _GEN_13;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_6_im <= 64'sh0; // @[Stap_Main.scala 128:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_6_im <= _GEN_12;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_7_re <= 64'sh0; // @[Stap_Main.scala 127:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_7_re <= _GEN_15;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_7_im <= 64'sh0; // @[Stap_Main.scala 128:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_7_im <= _GEN_14;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_8_re <= 64'sh0; // @[Stap_Main.scala 127:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_8_re <= _GEN_17;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_8_im <= 64'sh0; // @[Stap_Main.scala 128:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_8_im <= _GEN_16;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_9_re <= 64'sh0; // @[Stap_Main.scala 127:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_9_re <= _GEN_19;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_9_im <= 64'sh0; // @[Stap_Main.scala 128:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_9_im <= _GEN_18;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_10_re <= 64'sh0; // @[Stap_Main.scala 127:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_10_re <= _GEN_21;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_10_im <= 64'sh0; // @[Stap_Main.scala 128:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_10_im <= _GEN_20;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_11_re <= 64'sh0; // @[Stap_Main.scala 127:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_11_re <= _GEN_23;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_11_im <= 64'sh0; // @[Stap_Main.scala 128:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_11_im <= _GEN_22;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_12_re <= 64'sh0; // @[Stap_Main.scala 127:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_12_re <= _GEN_25;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_12_im <= 64'sh0; // @[Stap_Main.scala 128:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_12_im <= _GEN_24;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_13_re <= 64'sh0; // @[Stap_Main.scala 127:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_13_re <= _GEN_27;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_13_im <= 64'sh0; // @[Stap_Main.scala 128:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_13_im <= _GEN_26;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_14_re <= 64'sh0; // @[Stap_Main.scala 127:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_14_re <= _GEN_29;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_14_im <= 64'sh0; // @[Stap_Main.scala 128:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_14_im <= _GEN_28;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_15_re <= 64'sh0; // @[Stap_Main.scala 127:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_15_re <= _GEN_31;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_15_im <= 64'sh0; // @[Stap_Main.scala 128:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (status == 8'h2) begin // @[Stap_Main.scala 147:32]
          matrix_R_15_im <= _GEN_30;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_0_re <= 64'sh0; // @[Stap_Main.scala 133:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_0_re <= _GEN_1007;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_0_im <= 64'sh0; // @[Stap_Main.scala 134:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_0_im <= _GEN_1006;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_1_re <= 64'sh0; // @[Stap_Main.scala 133:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_1_re <= _GEN_1009;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_1_im <= 64'sh0; // @[Stap_Main.scala 134:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_1_im <= _GEN_1008;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_2_re <= 64'sh0; // @[Stap_Main.scala 133:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_2_re <= _GEN_1011;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_2_im <= 64'sh0; // @[Stap_Main.scala 134:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_2_im <= _GEN_1010;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_3_re <= 64'sh0; // @[Stap_Main.scala 133:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_3_re <= _GEN_1013;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_3_im <= 64'sh0; // @[Stap_Main.scala 134:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_3_im <= _GEN_1012;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_4_re <= 64'sh0; // @[Stap_Main.scala 133:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_4_re <= _GEN_1015;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_4_im <= 64'sh0; // @[Stap_Main.scala 134:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_4_im <= _GEN_1014;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_5_re <= 64'sh0; // @[Stap_Main.scala 133:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_5_re <= _GEN_1017;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_5_im <= 64'sh0; // @[Stap_Main.scala 134:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_5_im <= _GEN_1016;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_6_re <= 64'sh0; // @[Stap_Main.scala 133:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_6_re <= _GEN_1019;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_6_im <= 64'sh0; // @[Stap_Main.scala 134:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_6_im <= _GEN_1018;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_7_re <= 64'sh0; // @[Stap_Main.scala 133:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_7_re <= _GEN_1021;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_7_im <= 64'sh0; // @[Stap_Main.scala 134:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_7_im <= _GEN_1020;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_8_re <= 64'sh0; // @[Stap_Main.scala 133:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_8_re <= _GEN_1023;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_8_im <= 64'sh0; // @[Stap_Main.scala 134:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_8_im <= _GEN_1022;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_9_re <= 64'sh0; // @[Stap_Main.scala 133:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_9_re <= _GEN_1025;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_L_9_im <= 64'sh0; // @[Stap_Main.scala 134:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_L_9_im <= _GEN_1024;
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_0_re <= _GEN_1048;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_0_im <= _GEN_1047;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_1_re <= _GEN_1050;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_1_im <= _GEN_1049;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_2_re <= _GEN_1052;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_2_im <= _GEN_1051;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_3_re <= _GEN_1054;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_3_im <= _GEN_1053;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_4_re <= _GEN_1056;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_4_im <= _GEN_1055;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_5_re <= _GEN_1058;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_5_im <= _GEN_1057;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_6_re <= _GEN_1060;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_6_im <= _GEN_1059;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_7_re <= _GEN_1062;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_7_im <= _GEN_1061;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_8_re <= _GEN_1064;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_8_im <= _GEN_1063;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_9_re <= _GEN_1066;
          end
        end
      end
    end
    if (!(io_reset)) begin // @[Stap_Main.scala 114:18]
      if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
        if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
          if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
            matrix_L_inv_9_im <= _GEN_1065;
          end
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_0_re <= 64'sh0; // @[Stap_Main.scala 129:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_0_re <= _GEN_1133;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_0_im <= 64'sh0; // @[Stap_Main.scala 130:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_0_im <= _GEN_1132;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_1_re <= 64'sh0; // @[Stap_Main.scala 129:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_1_re <= _GEN_1135;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_1_im <= 64'sh0; // @[Stap_Main.scala 130:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_1_im <= _GEN_1134;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_2_re <= 64'sh0; // @[Stap_Main.scala 129:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_2_re <= _GEN_1137;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_2_im <= 64'sh0; // @[Stap_Main.scala 130:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_2_im <= _GEN_1136;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_3_re <= 64'sh0; // @[Stap_Main.scala 129:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_3_re <= _GEN_1139;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_3_im <= 64'sh0; // @[Stap_Main.scala 130:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_3_im <= _GEN_1138;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_4_re <= 64'sh0; // @[Stap_Main.scala 129:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_4_re <= _GEN_1141;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_4_im <= 64'sh0; // @[Stap_Main.scala 130:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_4_im <= _GEN_1140;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_5_re <= 64'sh0; // @[Stap_Main.scala 129:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_5_re <= _GEN_1143;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_5_im <= 64'sh0; // @[Stap_Main.scala 130:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_5_im <= _GEN_1142;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_6_re <= 64'sh0; // @[Stap_Main.scala 129:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_6_re <= _GEN_1145;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_6_im <= 64'sh0; // @[Stap_Main.scala 130:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_6_im <= _GEN_1144;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_7_re <= 64'sh0; // @[Stap_Main.scala 129:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_7_re <= _GEN_1147;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_7_im <= 64'sh0; // @[Stap_Main.scala 130:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_7_im <= _GEN_1146;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_8_re <= 64'sh0; // @[Stap_Main.scala 129:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_8_re <= _GEN_1149;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_8_im <= 64'sh0; // @[Stap_Main.scala 130:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_8_im <= _GEN_1148;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_9_re <= 64'sh0; // @[Stap_Main.scala 129:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_9_re <= _GEN_1151;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_9_im <= 64'sh0; // @[Stap_Main.scala 130:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_9_im <= _GEN_1150;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_10_re <= 64'sh0; // @[Stap_Main.scala 129:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_10_re <= _GEN_1153;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_10_im <= 64'sh0; // @[Stap_Main.scala 130:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_10_im <= _GEN_1152;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_11_re <= 64'sh0; // @[Stap_Main.scala 129:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_11_re <= _GEN_1155;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_11_im <= 64'sh0; // @[Stap_Main.scala 130:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_11_im <= _GEN_1154;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_12_re <= 64'sh0; // @[Stap_Main.scala 129:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_12_re <= _GEN_1157;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_12_im <= 64'sh0; // @[Stap_Main.scala 130:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_12_im <= _GEN_1156;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_13_re <= 64'sh0; // @[Stap_Main.scala 129:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_13_re <= _GEN_1159;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_13_im <= 64'sh0; // @[Stap_Main.scala 130:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_13_im <= _GEN_1158;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_14_re <= 64'sh0; // @[Stap_Main.scala 129:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_14_re <= _GEN_1161;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_14_im <= 64'sh0; // @[Stap_Main.scala 130:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_14_im <= _GEN_1160;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_15_re <= 64'sh0; // @[Stap_Main.scala 129:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_15_re <= _GEN_1163;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_R_inv_15_im <= 64'sh0; // @[Stap_Main.scala 130:26]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_R_inv_15_im <= _GEN_1162;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_w_0_re <= 64'sh0; // @[Stap_Main.scala 123:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_w_0_re <= _GEN_1206;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_w_0_im <= 64'sh0; // @[Stap_Main.scala 124:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_w_0_im <= _GEN_1205;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_w_1_re <= 64'sh0; // @[Stap_Main.scala 123:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_w_1_re <= _GEN_1208;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_w_1_im <= 64'sh0; // @[Stap_Main.scala 124:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_w_1_im <= _GEN_1207;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_w_2_re <= 64'sh0; // @[Stap_Main.scala 123:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_w_2_re <= _GEN_1210;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_w_2_im <= 64'sh0; // @[Stap_Main.scala 124:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_w_2_im <= _GEN_1209;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_w_3_re <= 64'sh0; // @[Stap_Main.scala 123:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_w_3_re <= _GEN_1212;
        end
      end
    end
    if (io_reset) begin // @[Stap_Main.scala 114:18]
      matrix_w_3_im <= 64'sh0; // @[Stap_Main.scala 124:22]
    end else if (!(io_ready)) begin // @[Stap_Main.scala 137:24]
      if (!(status == 8'h1)) begin // @[Stap_Main.scala 142:26]
        if (!(status == 8'h2)) begin // @[Stap_Main.scala 147:32]
          matrix_w_3_im <= _GEN_1211;
        end
      end
    end
    if (reset) begin // @[Stap_Main.scala 66:29]
      status <= 8'h0; // @[Stap_Main.scala 66:29]
    end else if (io_reset) begin // @[Stap_Main.scala 114:18]
      status <= 8'h0; // @[Stap_Main.scala 136:12]
    end else if (io_ready) begin // @[Stap_Main.scala 137:24]
      status <= 8'h1; // @[Stap_Main.scala 140:12]
    end else if (status == 8'h1) begin // @[Stap_Main.scala 142:26]
      status <= _status_T_1; // @[Stap_Main.scala 146:14]
    end else begin
      status <= _GEN_1246;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  matrix_x_in_0_re = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  matrix_x_in_0_im = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  matrix_x_in_1_re = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  matrix_x_in_1_im = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  matrix_x_in_2_re = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  matrix_x_in_2_im = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  matrix_x_in_3_re = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  matrix_x_in_3_im = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  matrix_x_in_4_re = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  matrix_x_in_4_im = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  matrix_x_in_5_re = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  matrix_x_in_5_im = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  matrix_x_in_6_re = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  matrix_x_in_6_im = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  matrix_x_in_7_re = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  matrix_x_in_7_im = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  matrix_S_0_re = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  matrix_S_0_im = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  matrix_S_1_re = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  matrix_S_1_im = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  matrix_S_2_re = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  matrix_S_2_im = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  matrix_S_3_re = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  matrix_S_3_im = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  matrix_R_0_re = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  matrix_R_0_im = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  matrix_R_1_re = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  matrix_R_1_im = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  matrix_R_2_re = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  matrix_R_2_im = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  matrix_R_3_re = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  matrix_R_3_im = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  matrix_R_4_re = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  matrix_R_4_im = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  matrix_R_5_re = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  matrix_R_5_im = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  matrix_R_6_re = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  matrix_R_6_im = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  matrix_R_7_re = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  matrix_R_7_im = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  matrix_R_8_re = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  matrix_R_8_im = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  matrix_R_9_re = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  matrix_R_9_im = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  matrix_R_10_re = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  matrix_R_10_im = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  matrix_R_11_re = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  matrix_R_11_im = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  matrix_R_12_re = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  matrix_R_12_im = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  matrix_R_13_re = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  matrix_R_13_im = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  matrix_R_14_re = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  matrix_R_14_im = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  matrix_R_15_re = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  matrix_R_15_im = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  matrix_L_0_re = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  matrix_L_0_im = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  matrix_L_1_re = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  matrix_L_1_im = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  matrix_L_2_re = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  matrix_L_2_im = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  matrix_L_3_re = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  matrix_L_3_im = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  matrix_L_4_re = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  matrix_L_4_im = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  matrix_L_5_re = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  matrix_L_5_im = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  matrix_L_6_re = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  matrix_L_6_im = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  matrix_L_7_re = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  matrix_L_7_im = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  matrix_L_8_re = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  matrix_L_8_im = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  matrix_L_9_re = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  matrix_L_9_im = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  matrix_L_inv_0_re = _RAND_76[63:0];
  _RAND_77 = {2{`RANDOM}};
  matrix_L_inv_0_im = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  matrix_L_inv_1_re = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  matrix_L_inv_1_im = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  matrix_L_inv_2_re = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  matrix_L_inv_2_im = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  matrix_L_inv_3_re = _RAND_82[63:0];
  _RAND_83 = {2{`RANDOM}};
  matrix_L_inv_3_im = _RAND_83[63:0];
  _RAND_84 = {2{`RANDOM}};
  matrix_L_inv_4_re = _RAND_84[63:0];
  _RAND_85 = {2{`RANDOM}};
  matrix_L_inv_4_im = _RAND_85[63:0];
  _RAND_86 = {2{`RANDOM}};
  matrix_L_inv_5_re = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  matrix_L_inv_5_im = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  matrix_L_inv_6_re = _RAND_88[63:0];
  _RAND_89 = {2{`RANDOM}};
  matrix_L_inv_6_im = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  matrix_L_inv_7_re = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  matrix_L_inv_7_im = _RAND_91[63:0];
  _RAND_92 = {2{`RANDOM}};
  matrix_L_inv_8_re = _RAND_92[63:0];
  _RAND_93 = {2{`RANDOM}};
  matrix_L_inv_8_im = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  matrix_L_inv_9_re = _RAND_94[63:0];
  _RAND_95 = {2{`RANDOM}};
  matrix_L_inv_9_im = _RAND_95[63:0];
  _RAND_96 = {2{`RANDOM}};
  matrix_R_inv_0_re = _RAND_96[63:0];
  _RAND_97 = {2{`RANDOM}};
  matrix_R_inv_0_im = _RAND_97[63:0];
  _RAND_98 = {2{`RANDOM}};
  matrix_R_inv_1_re = _RAND_98[63:0];
  _RAND_99 = {2{`RANDOM}};
  matrix_R_inv_1_im = _RAND_99[63:0];
  _RAND_100 = {2{`RANDOM}};
  matrix_R_inv_2_re = _RAND_100[63:0];
  _RAND_101 = {2{`RANDOM}};
  matrix_R_inv_2_im = _RAND_101[63:0];
  _RAND_102 = {2{`RANDOM}};
  matrix_R_inv_3_re = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  matrix_R_inv_3_im = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  matrix_R_inv_4_re = _RAND_104[63:0];
  _RAND_105 = {2{`RANDOM}};
  matrix_R_inv_4_im = _RAND_105[63:0];
  _RAND_106 = {2{`RANDOM}};
  matrix_R_inv_5_re = _RAND_106[63:0];
  _RAND_107 = {2{`RANDOM}};
  matrix_R_inv_5_im = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  matrix_R_inv_6_re = _RAND_108[63:0];
  _RAND_109 = {2{`RANDOM}};
  matrix_R_inv_6_im = _RAND_109[63:0];
  _RAND_110 = {2{`RANDOM}};
  matrix_R_inv_7_re = _RAND_110[63:0];
  _RAND_111 = {2{`RANDOM}};
  matrix_R_inv_7_im = _RAND_111[63:0];
  _RAND_112 = {2{`RANDOM}};
  matrix_R_inv_8_re = _RAND_112[63:0];
  _RAND_113 = {2{`RANDOM}};
  matrix_R_inv_8_im = _RAND_113[63:0];
  _RAND_114 = {2{`RANDOM}};
  matrix_R_inv_9_re = _RAND_114[63:0];
  _RAND_115 = {2{`RANDOM}};
  matrix_R_inv_9_im = _RAND_115[63:0];
  _RAND_116 = {2{`RANDOM}};
  matrix_R_inv_10_re = _RAND_116[63:0];
  _RAND_117 = {2{`RANDOM}};
  matrix_R_inv_10_im = _RAND_117[63:0];
  _RAND_118 = {2{`RANDOM}};
  matrix_R_inv_11_re = _RAND_118[63:0];
  _RAND_119 = {2{`RANDOM}};
  matrix_R_inv_11_im = _RAND_119[63:0];
  _RAND_120 = {2{`RANDOM}};
  matrix_R_inv_12_re = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  matrix_R_inv_12_im = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  matrix_R_inv_13_re = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  matrix_R_inv_13_im = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  matrix_R_inv_14_re = _RAND_124[63:0];
  _RAND_125 = {2{`RANDOM}};
  matrix_R_inv_14_im = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  matrix_R_inv_15_re = _RAND_126[63:0];
  _RAND_127 = {2{`RANDOM}};
  matrix_R_inv_15_im = _RAND_127[63:0];
  _RAND_128 = {2{`RANDOM}};
  matrix_w_0_re = _RAND_128[63:0];
  _RAND_129 = {2{`RANDOM}};
  matrix_w_0_im = _RAND_129[63:0];
  _RAND_130 = {2{`RANDOM}};
  matrix_w_1_re = _RAND_130[63:0];
  _RAND_131 = {2{`RANDOM}};
  matrix_w_1_im = _RAND_131[63:0];
  _RAND_132 = {2{`RANDOM}};
  matrix_w_2_re = _RAND_132[63:0];
  _RAND_133 = {2{`RANDOM}};
  matrix_w_2_im = _RAND_133[63:0];
  _RAND_134 = {2{`RANDOM}};
  matrix_w_3_re = _RAND_134[63:0];
  _RAND_135 = {2{`RANDOM}};
  matrix_w_3_im = _RAND_135[63:0];
  _RAND_136 = {1{`RANDOM}};
  status = _RAND_136[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
