module ComplexMul(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  wire [31:0] _k1_T_2 = $signed(io_op1_re) + $signed(io_op1_im); // @[Complex_Operater.scala 38:35]
  wire [63:0] k1 = $signed(io_op2_re) * $signed(_k1_T_2); // @[Complex_Operater.scala 38:22]
  wire [31:0] _k2_T_2 = $signed(io_op2_im) - $signed(io_op2_re); // @[Complex_Operater.scala 39:35]
  wire [63:0] k2 = $signed(io_op1_re) * $signed(_k2_T_2); // @[Complex_Operater.scala 39:22]
  wire [31:0] _k3_T_2 = $signed(io_op2_re) + $signed(io_op2_im); // @[Complex_Operater.scala 40:35]
  wire [63:0] k3 = $signed(io_op1_im) * $signed(_k3_T_2); // @[Complex_Operater.scala 40:22]
  wire [63:0] _io_res_re_T_2 = $signed(k1) - $signed(k3); // @[Complex_Operater.scala 41:19]
  wire [63:0] _io_res_im_T_2 = $signed(k1) + $signed(k2); // @[Complex_Operater.scala 42:19]
  wire [43:0] _GEN_0 = _io_res_re_T_2[63:20]; // @[Complex_Operater.scala 41:13]
  wire [43:0] _GEN_2 = _io_res_im_T_2[63:20]; // @[Complex_Operater.scala 42:13]
  assign io_res_re = _GEN_0[31:0]; // @[Complex_Operater.scala 41:13]
  assign io_res_im = _GEN_2[31:0]; // @[Complex_Operater.scala 42:13]
endmodule
module ComplexAdd(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) + $signed(io_op2_re); // @[Complex_Operater.scala 7:26]
  assign io_res_im = $signed(io_op1_im) + $signed(io_op2_im); // @[Complex_Operater.scala 8:26]
endmodule
module PE(
  input         clock,
  input         io_reset,
  input  [31:0] io_in_x_re,
  input  [31:0] io_in_x_im,
  input  [31:0] io_in_y_re,
  input  [31:0] io_in_y_im,
  output [31:0] io_out_pe_re,
  output [31:0] io_out_pe_im,
  output [31:0] io_out_x_re,
  output [31:0] io_out_x_im,
  output [31:0] io_out_y_re,
  output [31:0] io_out_y_im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] pe_reg_mul_io_op1_re; // @[Complex_Operater.scala 47:21]
  wire [31:0] pe_reg_mul_io_op1_im; // @[Complex_Operater.scala 47:21]
  wire [31:0] pe_reg_mul_io_op2_re; // @[Complex_Operater.scala 47:21]
  wire [31:0] pe_reg_mul_io_op2_im; // @[Complex_Operater.scala 47:21]
  wire [31:0] pe_reg_mul_io_res_re; // @[Complex_Operater.scala 47:21]
  wire [31:0] pe_reg_mul_io_res_im; // @[Complex_Operater.scala 47:21]
  wire [31:0] pe_reg_add_io_op1_re; // @[Complex_Operater.scala 13:21]
  wire [31:0] pe_reg_add_io_op1_im; // @[Complex_Operater.scala 13:21]
  wire [31:0] pe_reg_add_io_op2_re; // @[Complex_Operater.scala 13:21]
  wire [31:0] pe_reg_add_io_op2_im; // @[Complex_Operater.scala 13:21]
  wire [31:0] pe_reg_add_io_res_re; // @[Complex_Operater.scala 13:21]
  wire [31:0] pe_reg_add_io_res_im; // @[Complex_Operater.scala 13:21]
  reg [31:0] pe_reg_re; // @[Matrix_Mul_V1.scala 29:28]
  reg [31:0] pe_reg_im; // @[Matrix_Mul_V1.scala 29:28]
  reg [31:0] x_reg_re; // @[Matrix_Mul_V1.scala 30:27]
  reg [31:0] x_reg_im; // @[Matrix_Mul_V1.scala 30:27]
  reg [31:0] y_reg_re; // @[Matrix_Mul_V1.scala 31:27]
  reg [31:0] y_reg_im; // @[Matrix_Mul_V1.scala 31:27]
  ComplexMul pe_reg_mul ( // @[Complex_Operater.scala 47:21]
    .io_op1_re(pe_reg_mul_io_op1_re),
    .io_op1_im(pe_reg_mul_io_op1_im),
    .io_op2_re(pe_reg_mul_io_op2_re),
    .io_op2_im(pe_reg_mul_io_op2_im),
    .io_res_re(pe_reg_mul_io_res_re),
    .io_res_im(pe_reg_mul_io_res_im)
  );
  ComplexAdd pe_reg_add ( // @[Complex_Operater.scala 13:21]
    .io_op1_re(pe_reg_add_io_op1_re),
    .io_op1_im(pe_reg_add_io_op1_im),
    .io_op2_re(pe_reg_add_io_op2_re),
    .io_op2_im(pe_reg_add_io_op2_im),
    .io_res_re(pe_reg_add_io_res_re),
    .io_res_im(pe_reg_add_io_res_im)
  );
  assign io_out_pe_re = pe_reg_re; // @[Matrix_Mul_V1.scala 50:13]
  assign io_out_pe_im = pe_reg_im; // @[Matrix_Mul_V1.scala 50:13]
  assign io_out_x_re = x_reg_re; // @[Matrix_Mul_V1.scala 51:12]
  assign io_out_x_im = x_reg_im; // @[Matrix_Mul_V1.scala 51:12]
  assign io_out_y_re = y_reg_re; // @[Matrix_Mul_V1.scala 52:12]
  assign io_out_y_im = y_reg_im; // @[Matrix_Mul_V1.scala 52:12]
  assign pe_reg_mul_io_op1_re = io_in_x_re; // @[Complex_Operater.scala 48:16]
  assign pe_reg_mul_io_op1_im = io_in_x_im; // @[Complex_Operater.scala 48:16]
  assign pe_reg_mul_io_op2_re = io_in_y_re; // @[Complex_Operater.scala 49:16]
  assign pe_reg_mul_io_op2_im = io_in_y_im; // @[Complex_Operater.scala 49:16]
  assign pe_reg_add_io_op1_re = pe_reg_re; // @[Complex_Operater.scala 14:16]
  assign pe_reg_add_io_op1_im = pe_reg_im; // @[Complex_Operater.scala 14:16]
  assign pe_reg_add_io_op2_re = pe_reg_mul_io_res_re; // @[Complex_Operater.scala 15:16]
  assign pe_reg_add_io_op2_im = pe_reg_mul_io_res_im; // @[Complex_Operater.scala 15:16]
  always @(posedge clock) begin
    if (io_reset) begin // @[Matrix_Mul_V1.scala 33:18]
      pe_reg_re <= 32'sh0; // @[Matrix_Mul_V1.scala 35:15]
    end else begin
      pe_reg_re <= pe_reg_add_io_res_re; // @[Matrix_Mul_V1.scala 43:12]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 33:18]
      pe_reg_im <= 32'sh0; // @[Matrix_Mul_V1.scala 36:15]
    end else begin
      pe_reg_im <= pe_reg_add_io_res_im; // @[Matrix_Mul_V1.scala 43:12]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 33:18]
      x_reg_re <= 32'sh0; // @[Matrix_Mul_V1.scala 37:14]
    end else begin
      x_reg_re <= io_in_x_re; // @[Matrix_Mul_V1.scala 45:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 33:18]
      x_reg_im <= 32'sh0; // @[Matrix_Mul_V1.scala 38:14]
    end else begin
      x_reg_im <= io_in_x_im; // @[Matrix_Mul_V1.scala 45:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 33:18]
      y_reg_re <= 32'sh0; // @[Matrix_Mul_V1.scala 39:14]
    end else begin
      y_reg_re <= io_in_y_re; // @[Matrix_Mul_V1.scala 46:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 33:18]
      y_reg_im <= 32'sh0; // @[Matrix_Mul_V1.scala 40:14]
    end else begin
      y_reg_im <= io_in_y_im; // @[Matrix_Mul_V1.scala 46:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pe_reg_re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  pe_reg_im = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  x_reg_re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  x_reg_im = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  y_reg_re = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  y_reg_im = _RAND_5[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module matrix_mul_v1(
  input         clock,
  input         reset,
  input         io_reset,
  input         io_ready,
  input  [31:0] io_matrixA_0_re,
  input  [31:0] io_matrixA_0_im,
  input  [31:0] io_matrixA_1_re,
  input  [31:0] io_matrixA_1_im,
  input  [31:0] io_matrixA_2_re,
  input  [31:0] io_matrixA_2_im,
  input  [31:0] io_matrixA_3_re,
  input  [31:0] io_matrixA_3_im,
  input  [31:0] io_matrixA_4_re,
  input  [31:0] io_matrixA_4_im,
  input  [31:0] io_matrixA_5_re,
  input  [31:0] io_matrixA_5_im,
  input  [31:0] io_matrixA_6_re,
  input  [31:0] io_matrixA_6_im,
  input  [31:0] io_matrixA_7_re,
  input  [31:0] io_matrixA_7_im,
  input  [31:0] io_matrixA_8_re,
  input  [31:0] io_matrixA_8_im,
  input  [31:0] io_matrixA_9_re,
  input  [31:0] io_matrixA_9_im,
  input  [31:0] io_matrixA_10_re,
  input  [31:0] io_matrixA_10_im,
  input  [31:0] io_matrixA_11_re,
  input  [31:0] io_matrixA_11_im,
  input  [31:0] io_matrixA_12_re,
  input  [31:0] io_matrixA_12_im,
  input  [31:0] io_matrixA_13_re,
  input  [31:0] io_matrixA_13_im,
  input  [31:0] io_matrixA_14_re,
  input  [31:0] io_matrixA_14_im,
  input  [31:0] io_matrixA_15_re,
  input  [31:0] io_matrixA_15_im,
  input  [31:0] io_matrixA_16_re,
  input  [31:0] io_matrixA_16_im,
  input  [31:0] io_matrixA_17_re,
  input  [31:0] io_matrixA_17_im,
  input  [31:0] io_matrixA_18_re,
  input  [31:0] io_matrixA_18_im,
  input  [31:0] io_matrixA_19_re,
  input  [31:0] io_matrixA_19_im,
  input  [31:0] io_matrixA_20_re,
  input  [31:0] io_matrixA_20_im,
  input  [31:0] io_matrixA_21_re,
  input  [31:0] io_matrixA_21_im,
  input  [31:0] io_matrixA_22_re,
  input  [31:0] io_matrixA_22_im,
  input  [31:0] io_matrixA_23_re,
  input  [31:0] io_matrixA_23_im,
  input  [31:0] io_matrixA_24_re,
  input  [31:0] io_matrixA_24_im,
  input  [31:0] io_matrixA_25_re,
  input  [31:0] io_matrixA_25_im,
  input  [31:0] io_matrixA_26_re,
  input  [31:0] io_matrixA_26_im,
  input  [31:0] io_matrixA_27_re,
  input  [31:0] io_matrixA_27_im,
  input  [31:0] io_matrixA_28_re,
  input  [31:0] io_matrixA_28_im,
  input  [31:0] io_matrixA_29_re,
  input  [31:0] io_matrixA_29_im,
  input  [31:0] io_matrixA_30_re,
  input  [31:0] io_matrixA_30_im,
  input  [31:0] io_matrixA_31_re,
  input  [31:0] io_matrixA_31_im,
  input  [31:0] io_matrixA_32_re,
  input  [31:0] io_matrixA_32_im,
  input  [31:0] io_matrixA_33_re,
  input  [31:0] io_matrixA_33_im,
  input  [31:0] io_matrixA_34_re,
  input  [31:0] io_matrixA_34_im,
  input  [31:0] io_matrixA_35_re,
  input  [31:0] io_matrixA_35_im,
  input  [31:0] io_matrixA_36_re,
  input  [31:0] io_matrixA_36_im,
  input  [31:0] io_matrixA_37_re,
  input  [31:0] io_matrixA_37_im,
  input  [31:0] io_matrixA_38_re,
  input  [31:0] io_matrixA_38_im,
  input  [31:0] io_matrixA_39_re,
  input  [31:0] io_matrixA_39_im,
  input  [31:0] io_matrixA_40_re,
  input  [31:0] io_matrixA_40_im,
  input  [31:0] io_matrixA_41_re,
  input  [31:0] io_matrixA_41_im,
  input  [31:0] io_matrixA_42_re,
  input  [31:0] io_matrixA_42_im,
  input  [31:0] io_matrixA_43_re,
  input  [31:0] io_matrixA_43_im,
  input  [31:0] io_matrixA_44_re,
  input  [31:0] io_matrixA_44_im,
  input  [31:0] io_matrixA_45_re,
  input  [31:0] io_matrixA_45_im,
  input  [31:0] io_matrixA_46_re,
  input  [31:0] io_matrixA_46_im,
  input  [31:0] io_matrixA_47_re,
  input  [31:0] io_matrixA_47_im,
  input  [31:0] io_matrixA_48_re,
  input  [31:0] io_matrixA_48_im,
  input  [31:0] io_matrixA_49_re,
  input  [31:0] io_matrixA_49_im,
  input  [31:0] io_matrixA_50_re,
  input  [31:0] io_matrixA_50_im,
  input  [31:0] io_matrixA_51_re,
  input  [31:0] io_matrixA_51_im,
  input  [31:0] io_matrixA_52_re,
  input  [31:0] io_matrixA_52_im,
  input  [31:0] io_matrixA_53_re,
  input  [31:0] io_matrixA_53_im,
  input  [31:0] io_matrixA_54_re,
  input  [31:0] io_matrixA_54_im,
  input  [31:0] io_matrixA_55_re,
  input  [31:0] io_matrixA_55_im,
  input  [31:0] io_matrixA_56_re,
  input  [31:0] io_matrixA_56_im,
  input  [31:0] io_matrixA_57_re,
  input  [31:0] io_matrixA_57_im,
  input  [31:0] io_matrixA_58_re,
  input  [31:0] io_matrixA_58_im,
  input  [31:0] io_matrixA_59_re,
  input  [31:0] io_matrixA_59_im,
  input  [31:0] io_matrixA_60_re,
  input  [31:0] io_matrixA_60_im,
  input  [31:0] io_matrixA_61_re,
  input  [31:0] io_matrixA_61_im,
  input  [31:0] io_matrixA_62_re,
  input  [31:0] io_matrixA_62_im,
  input  [31:0] io_matrixA_63_re,
  input  [31:0] io_matrixA_63_im,
  input  [31:0] io_matrixA_64_re,
  input  [31:0] io_matrixA_64_im,
  input  [31:0] io_matrixA_65_re,
  input  [31:0] io_matrixA_65_im,
  input  [31:0] io_matrixA_66_re,
  input  [31:0] io_matrixA_66_im,
  input  [31:0] io_matrixA_67_re,
  input  [31:0] io_matrixA_67_im,
  input  [31:0] io_matrixA_68_re,
  input  [31:0] io_matrixA_68_im,
  input  [31:0] io_matrixA_69_re,
  input  [31:0] io_matrixA_69_im,
  input  [31:0] io_matrixA_70_re,
  input  [31:0] io_matrixA_70_im,
  input  [31:0] io_matrixA_71_re,
  input  [31:0] io_matrixA_71_im,
  input  [31:0] io_matrixA_72_re,
  input  [31:0] io_matrixA_72_im,
  input  [31:0] io_matrixA_73_re,
  input  [31:0] io_matrixA_73_im,
  input  [31:0] io_matrixA_74_re,
  input  [31:0] io_matrixA_74_im,
  input  [31:0] io_matrixA_75_re,
  input  [31:0] io_matrixA_75_im,
  input  [31:0] io_matrixA_76_re,
  input  [31:0] io_matrixA_76_im,
  input  [31:0] io_matrixA_77_re,
  input  [31:0] io_matrixA_77_im,
  input  [31:0] io_matrixA_78_re,
  input  [31:0] io_matrixA_78_im,
  input  [31:0] io_matrixA_79_re,
  input  [31:0] io_matrixA_79_im,
  input  [31:0] io_matrixA_80_re,
  input  [31:0] io_matrixA_80_im,
  input  [31:0] io_matrixA_81_re,
  input  [31:0] io_matrixA_81_im,
  input  [31:0] io_matrixA_82_re,
  input  [31:0] io_matrixA_82_im,
  input  [31:0] io_matrixA_83_re,
  input  [31:0] io_matrixA_83_im,
  input  [31:0] io_matrixA_84_re,
  input  [31:0] io_matrixA_84_im,
  input  [31:0] io_matrixA_85_re,
  input  [31:0] io_matrixA_85_im,
  input  [31:0] io_matrixA_86_re,
  input  [31:0] io_matrixA_86_im,
  input  [31:0] io_matrixA_87_re,
  input  [31:0] io_matrixA_87_im,
  input  [31:0] io_matrixA_88_re,
  input  [31:0] io_matrixA_88_im,
  input  [31:0] io_matrixA_89_re,
  input  [31:0] io_matrixA_89_im,
  input  [31:0] io_matrixA_90_re,
  input  [31:0] io_matrixA_90_im,
  input  [31:0] io_matrixA_91_re,
  input  [31:0] io_matrixA_91_im,
  input  [31:0] io_matrixA_92_re,
  input  [31:0] io_matrixA_92_im,
  input  [31:0] io_matrixA_93_re,
  input  [31:0] io_matrixA_93_im,
  input  [31:0] io_matrixA_94_re,
  input  [31:0] io_matrixA_94_im,
  input  [31:0] io_matrixA_95_re,
  input  [31:0] io_matrixA_95_im,
  input  [31:0] io_matrixA_96_re,
  input  [31:0] io_matrixA_96_im,
  input  [31:0] io_matrixA_97_re,
  input  [31:0] io_matrixA_97_im,
  input  [31:0] io_matrixA_98_re,
  input  [31:0] io_matrixA_98_im,
  input  [31:0] io_matrixA_99_re,
  input  [31:0] io_matrixA_99_im,
  input  [31:0] io_matrixB_0_re,
  input  [31:0] io_matrixB_0_im,
  input  [31:0] io_matrixB_1_re,
  input  [31:0] io_matrixB_1_im,
  input  [31:0] io_matrixB_2_re,
  input  [31:0] io_matrixB_2_im,
  input  [31:0] io_matrixB_3_re,
  input  [31:0] io_matrixB_3_im,
  input  [31:0] io_matrixB_4_re,
  input  [31:0] io_matrixB_4_im,
  input  [31:0] io_matrixB_5_re,
  input  [31:0] io_matrixB_5_im,
  input  [31:0] io_matrixB_6_re,
  input  [31:0] io_matrixB_6_im,
  input  [31:0] io_matrixB_7_re,
  input  [31:0] io_matrixB_7_im,
  input  [31:0] io_matrixB_8_re,
  input  [31:0] io_matrixB_8_im,
  input  [31:0] io_matrixB_9_re,
  input  [31:0] io_matrixB_9_im,
  input  [31:0] io_matrixB_10_re,
  input  [31:0] io_matrixB_10_im,
  input  [31:0] io_matrixB_11_re,
  input  [31:0] io_matrixB_11_im,
  input  [31:0] io_matrixB_12_re,
  input  [31:0] io_matrixB_12_im,
  input  [31:0] io_matrixB_13_re,
  input  [31:0] io_matrixB_13_im,
  input  [31:0] io_matrixB_14_re,
  input  [31:0] io_matrixB_14_im,
  input  [31:0] io_matrixB_15_re,
  input  [31:0] io_matrixB_15_im,
  input  [31:0] io_matrixB_16_re,
  input  [31:0] io_matrixB_16_im,
  input  [31:0] io_matrixB_17_re,
  input  [31:0] io_matrixB_17_im,
  input  [31:0] io_matrixB_18_re,
  input  [31:0] io_matrixB_18_im,
  input  [31:0] io_matrixB_19_re,
  input  [31:0] io_matrixB_19_im,
  input  [31:0] io_matrixB_20_re,
  input  [31:0] io_matrixB_20_im,
  input  [31:0] io_matrixB_21_re,
  input  [31:0] io_matrixB_21_im,
  input  [31:0] io_matrixB_22_re,
  input  [31:0] io_matrixB_22_im,
  input  [31:0] io_matrixB_23_re,
  input  [31:0] io_matrixB_23_im,
  input  [31:0] io_matrixB_24_re,
  input  [31:0] io_matrixB_24_im,
  input  [31:0] io_matrixB_25_re,
  input  [31:0] io_matrixB_25_im,
  input  [31:0] io_matrixB_26_re,
  input  [31:0] io_matrixB_26_im,
  input  [31:0] io_matrixB_27_re,
  input  [31:0] io_matrixB_27_im,
  input  [31:0] io_matrixB_28_re,
  input  [31:0] io_matrixB_28_im,
  input  [31:0] io_matrixB_29_re,
  input  [31:0] io_matrixB_29_im,
  input  [31:0] io_matrixB_30_re,
  input  [31:0] io_matrixB_30_im,
  input  [31:0] io_matrixB_31_re,
  input  [31:0] io_matrixB_31_im,
  input  [31:0] io_matrixB_32_re,
  input  [31:0] io_matrixB_32_im,
  input  [31:0] io_matrixB_33_re,
  input  [31:0] io_matrixB_33_im,
  input  [31:0] io_matrixB_34_re,
  input  [31:0] io_matrixB_34_im,
  input  [31:0] io_matrixB_35_re,
  input  [31:0] io_matrixB_35_im,
  input  [31:0] io_matrixB_36_re,
  input  [31:0] io_matrixB_36_im,
  input  [31:0] io_matrixB_37_re,
  input  [31:0] io_matrixB_37_im,
  input  [31:0] io_matrixB_38_re,
  input  [31:0] io_matrixB_38_im,
  input  [31:0] io_matrixB_39_re,
  input  [31:0] io_matrixB_39_im,
  input  [31:0] io_matrixB_40_re,
  input  [31:0] io_matrixB_40_im,
  input  [31:0] io_matrixB_41_re,
  input  [31:0] io_matrixB_41_im,
  input  [31:0] io_matrixB_42_re,
  input  [31:0] io_matrixB_42_im,
  input  [31:0] io_matrixB_43_re,
  input  [31:0] io_matrixB_43_im,
  input  [31:0] io_matrixB_44_re,
  input  [31:0] io_matrixB_44_im,
  input  [31:0] io_matrixB_45_re,
  input  [31:0] io_matrixB_45_im,
  input  [31:0] io_matrixB_46_re,
  input  [31:0] io_matrixB_46_im,
  input  [31:0] io_matrixB_47_re,
  input  [31:0] io_matrixB_47_im,
  input  [31:0] io_matrixB_48_re,
  input  [31:0] io_matrixB_48_im,
  input  [31:0] io_matrixB_49_re,
  input  [31:0] io_matrixB_49_im,
  input  [31:0] io_matrixB_50_re,
  input  [31:0] io_matrixB_50_im,
  input  [31:0] io_matrixB_51_re,
  input  [31:0] io_matrixB_51_im,
  input  [31:0] io_matrixB_52_re,
  input  [31:0] io_matrixB_52_im,
  input  [31:0] io_matrixB_53_re,
  input  [31:0] io_matrixB_53_im,
  input  [31:0] io_matrixB_54_re,
  input  [31:0] io_matrixB_54_im,
  input  [31:0] io_matrixB_55_re,
  input  [31:0] io_matrixB_55_im,
  input  [31:0] io_matrixB_56_re,
  input  [31:0] io_matrixB_56_im,
  input  [31:0] io_matrixB_57_re,
  input  [31:0] io_matrixB_57_im,
  input  [31:0] io_matrixB_58_re,
  input  [31:0] io_matrixB_58_im,
  input  [31:0] io_matrixB_59_re,
  input  [31:0] io_matrixB_59_im,
  input  [31:0] io_matrixB_60_re,
  input  [31:0] io_matrixB_60_im,
  input  [31:0] io_matrixB_61_re,
  input  [31:0] io_matrixB_61_im,
  input  [31:0] io_matrixB_62_re,
  input  [31:0] io_matrixB_62_im,
  input  [31:0] io_matrixB_63_re,
  input  [31:0] io_matrixB_63_im,
  input  [31:0] io_matrixB_64_re,
  input  [31:0] io_matrixB_64_im,
  input  [31:0] io_matrixB_65_re,
  input  [31:0] io_matrixB_65_im,
  input  [31:0] io_matrixB_66_re,
  input  [31:0] io_matrixB_66_im,
  input  [31:0] io_matrixB_67_re,
  input  [31:0] io_matrixB_67_im,
  input  [31:0] io_matrixB_68_re,
  input  [31:0] io_matrixB_68_im,
  input  [31:0] io_matrixB_69_re,
  input  [31:0] io_matrixB_69_im,
  input  [31:0] io_matrixB_70_re,
  input  [31:0] io_matrixB_70_im,
  input  [31:0] io_matrixB_71_re,
  input  [31:0] io_matrixB_71_im,
  input  [31:0] io_matrixB_72_re,
  input  [31:0] io_matrixB_72_im,
  input  [31:0] io_matrixB_73_re,
  input  [31:0] io_matrixB_73_im,
  input  [31:0] io_matrixB_74_re,
  input  [31:0] io_matrixB_74_im,
  input  [31:0] io_matrixB_75_re,
  input  [31:0] io_matrixB_75_im,
  input  [31:0] io_matrixB_76_re,
  input  [31:0] io_matrixB_76_im,
  input  [31:0] io_matrixB_77_re,
  input  [31:0] io_matrixB_77_im,
  input  [31:0] io_matrixB_78_re,
  input  [31:0] io_matrixB_78_im,
  input  [31:0] io_matrixB_79_re,
  input  [31:0] io_matrixB_79_im,
  input  [31:0] io_matrixB_80_re,
  input  [31:0] io_matrixB_80_im,
  input  [31:0] io_matrixB_81_re,
  input  [31:0] io_matrixB_81_im,
  input  [31:0] io_matrixB_82_re,
  input  [31:0] io_matrixB_82_im,
  input  [31:0] io_matrixB_83_re,
  input  [31:0] io_matrixB_83_im,
  input  [31:0] io_matrixB_84_re,
  input  [31:0] io_matrixB_84_im,
  input  [31:0] io_matrixB_85_re,
  input  [31:0] io_matrixB_85_im,
  input  [31:0] io_matrixB_86_re,
  input  [31:0] io_matrixB_86_im,
  input  [31:0] io_matrixB_87_re,
  input  [31:0] io_matrixB_87_im,
  input  [31:0] io_matrixB_88_re,
  input  [31:0] io_matrixB_88_im,
  input  [31:0] io_matrixB_89_re,
  input  [31:0] io_matrixB_89_im,
  input  [31:0] io_matrixB_90_re,
  input  [31:0] io_matrixB_90_im,
  input  [31:0] io_matrixB_91_re,
  input  [31:0] io_matrixB_91_im,
  input  [31:0] io_matrixB_92_re,
  input  [31:0] io_matrixB_92_im,
  input  [31:0] io_matrixB_93_re,
  input  [31:0] io_matrixB_93_im,
  input  [31:0] io_matrixB_94_re,
  input  [31:0] io_matrixB_94_im,
  input  [31:0] io_matrixB_95_re,
  input  [31:0] io_matrixB_95_im,
  input  [31:0] io_matrixB_96_re,
  input  [31:0] io_matrixB_96_im,
  input  [31:0] io_matrixB_97_re,
  input  [31:0] io_matrixB_97_im,
  input  [31:0] io_matrixB_98_re,
  input  [31:0] io_matrixB_98_im,
  input  [31:0] io_matrixB_99_re,
  input  [31:0] io_matrixB_99_im,
  output [31:0] io_matrixC_0_re,
  output [31:0] io_matrixC_0_im,
  output [31:0] io_matrixC_1_re,
  output [31:0] io_matrixC_1_im,
  output [31:0] io_matrixC_2_re,
  output [31:0] io_matrixC_2_im,
  output [31:0] io_matrixC_3_re,
  output [31:0] io_matrixC_3_im,
  output [31:0] io_matrixC_4_re,
  output [31:0] io_matrixC_4_im,
  output [31:0] io_matrixC_5_re,
  output [31:0] io_matrixC_5_im,
  output [31:0] io_matrixC_6_re,
  output [31:0] io_matrixC_6_im,
  output [31:0] io_matrixC_7_re,
  output [31:0] io_matrixC_7_im,
  output [31:0] io_matrixC_8_re,
  output [31:0] io_matrixC_8_im,
  output [31:0] io_matrixC_9_re,
  output [31:0] io_matrixC_9_im,
  output [31:0] io_matrixC_10_re,
  output [31:0] io_matrixC_10_im,
  output [31:0] io_matrixC_11_re,
  output [31:0] io_matrixC_11_im,
  output [31:0] io_matrixC_12_re,
  output [31:0] io_matrixC_12_im,
  output [31:0] io_matrixC_13_re,
  output [31:0] io_matrixC_13_im,
  output [31:0] io_matrixC_14_re,
  output [31:0] io_matrixC_14_im,
  output [31:0] io_matrixC_15_re,
  output [31:0] io_matrixC_15_im,
  output [31:0] io_matrixC_16_re,
  output [31:0] io_matrixC_16_im,
  output [31:0] io_matrixC_17_re,
  output [31:0] io_matrixC_17_im,
  output [31:0] io_matrixC_18_re,
  output [31:0] io_matrixC_18_im,
  output [31:0] io_matrixC_19_re,
  output [31:0] io_matrixC_19_im,
  output [31:0] io_matrixC_20_re,
  output [31:0] io_matrixC_20_im,
  output [31:0] io_matrixC_21_re,
  output [31:0] io_matrixC_21_im,
  output [31:0] io_matrixC_22_re,
  output [31:0] io_matrixC_22_im,
  output [31:0] io_matrixC_23_re,
  output [31:0] io_matrixC_23_im,
  output [31:0] io_matrixC_24_re,
  output [31:0] io_matrixC_24_im,
  output [31:0] io_matrixC_25_re,
  output [31:0] io_matrixC_25_im,
  output [31:0] io_matrixC_26_re,
  output [31:0] io_matrixC_26_im,
  output [31:0] io_matrixC_27_re,
  output [31:0] io_matrixC_27_im,
  output [31:0] io_matrixC_28_re,
  output [31:0] io_matrixC_28_im,
  output [31:0] io_matrixC_29_re,
  output [31:0] io_matrixC_29_im,
  output [31:0] io_matrixC_30_re,
  output [31:0] io_matrixC_30_im,
  output [31:0] io_matrixC_31_re,
  output [31:0] io_matrixC_31_im,
  output [31:0] io_matrixC_32_re,
  output [31:0] io_matrixC_32_im,
  output [31:0] io_matrixC_33_re,
  output [31:0] io_matrixC_33_im,
  output [31:0] io_matrixC_34_re,
  output [31:0] io_matrixC_34_im,
  output [31:0] io_matrixC_35_re,
  output [31:0] io_matrixC_35_im,
  output [31:0] io_matrixC_36_re,
  output [31:0] io_matrixC_36_im,
  output [31:0] io_matrixC_37_re,
  output [31:0] io_matrixC_37_im,
  output [31:0] io_matrixC_38_re,
  output [31:0] io_matrixC_38_im,
  output [31:0] io_matrixC_39_re,
  output [31:0] io_matrixC_39_im,
  output [31:0] io_matrixC_40_re,
  output [31:0] io_matrixC_40_im,
  output [31:0] io_matrixC_41_re,
  output [31:0] io_matrixC_41_im,
  output [31:0] io_matrixC_42_re,
  output [31:0] io_matrixC_42_im,
  output [31:0] io_matrixC_43_re,
  output [31:0] io_matrixC_43_im,
  output [31:0] io_matrixC_44_re,
  output [31:0] io_matrixC_44_im,
  output [31:0] io_matrixC_45_re,
  output [31:0] io_matrixC_45_im,
  output [31:0] io_matrixC_46_re,
  output [31:0] io_matrixC_46_im,
  output [31:0] io_matrixC_47_re,
  output [31:0] io_matrixC_47_im,
  output [31:0] io_matrixC_48_re,
  output [31:0] io_matrixC_48_im,
  output [31:0] io_matrixC_49_re,
  output [31:0] io_matrixC_49_im,
  output [31:0] io_matrixC_50_re,
  output [31:0] io_matrixC_50_im,
  output [31:0] io_matrixC_51_re,
  output [31:0] io_matrixC_51_im,
  output [31:0] io_matrixC_52_re,
  output [31:0] io_matrixC_52_im,
  output [31:0] io_matrixC_53_re,
  output [31:0] io_matrixC_53_im,
  output [31:0] io_matrixC_54_re,
  output [31:0] io_matrixC_54_im,
  output [31:0] io_matrixC_55_re,
  output [31:0] io_matrixC_55_im,
  output [31:0] io_matrixC_56_re,
  output [31:0] io_matrixC_56_im,
  output [31:0] io_matrixC_57_re,
  output [31:0] io_matrixC_57_im,
  output [31:0] io_matrixC_58_re,
  output [31:0] io_matrixC_58_im,
  output [31:0] io_matrixC_59_re,
  output [31:0] io_matrixC_59_im,
  output [31:0] io_matrixC_60_re,
  output [31:0] io_matrixC_60_im,
  output [31:0] io_matrixC_61_re,
  output [31:0] io_matrixC_61_im,
  output [31:0] io_matrixC_62_re,
  output [31:0] io_matrixC_62_im,
  output [31:0] io_matrixC_63_re,
  output [31:0] io_matrixC_63_im,
  output [31:0] io_matrixC_64_re,
  output [31:0] io_matrixC_64_im,
  output [31:0] io_matrixC_65_re,
  output [31:0] io_matrixC_65_im,
  output [31:0] io_matrixC_66_re,
  output [31:0] io_matrixC_66_im,
  output [31:0] io_matrixC_67_re,
  output [31:0] io_matrixC_67_im,
  output [31:0] io_matrixC_68_re,
  output [31:0] io_matrixC_68_im,
  output [31:0] io_matrixC_69_re,
  output [31:0] io_matrixC_69_im,
  output [31:0] io_matrixC_70_re,
  output [31:0] io_matrixC_70_im,
  output [31:0] io_matrixC_71_re,
  output [31:0] io_matrixC_71_im,
  output [31:0] io_matrixC_72_re,
  output [31:0] io_matrixC_72_im,
  output [31:0] io_matrixC_73_re,
  output [31:0] io_matrixC_73_im,
  output [31:0] io_matrixC_74_re,
  output [31:0] io_matrixC_74_im,
  output [31:0] io_matrixC_75_re,
  output [31:0] io_matrixC_75_im,
  output [31:0] io_matrixC_76_re,
  output [31:0] io_matrixC_76_im,
  output [31:0] io_matrixC_77_re,
  output [31:0] io_matrixC_77_im,
  output [31:0] io_matrixC_78_re,
  output [31:0] io_matrixC_78_im,
  output [31:0] io_matrixC_79_re,
  output [31:0] io_matrixC_79_im,
  output [31:0] io_matrixC_80_re,
  output [31:0] io_matrixC_80_im,
  output [31:0] io_matrixC_81_re,
  output [31:0] io_matrixC_81_im,
  output [31:0] io_matrixC_82_re,
  output [31:0] io_matrixC_82_im,
  output [31:0] io_matrixC_83_re,
  output [31:0] io_matrixC_83_im,
  output [31:0] io_matrixC_84_re,
  output [31:0] io_matrixC_84_im,
  output [31:0] io_matrixC_85_re,
  output [31:0] io_matrixC_85_im,
  output [31:0] io_matrixC_86_re,
  output [31:0] io_matrixC_86_im,
  output [31:0] io_matrixC_87_re,
  output [31:0] io_matrixC_87_im,
  output [31:0] io_matrixC_88_re,
  output [31:0] io_matrixC_88_im,
  output [31:0] io_matrixC_89_re,
  output [31:0] io_matrixC_89_im,
  output [31:0] io_matrixC_90_re,
  output [31:0] io_matrixC_90_im,
  output [31:0] io_matrixC_91_re,
  output [31:0] io_matrixC_91_im,
  output [31:0] io_matrixC_92_re,
  output [31:0] io_matrixC_92_im,
  output [31:0] io_matrixC_93_re,
  output [31:0] io_matrixC_93_im,
  output [31:0] io_matrixC_94_re,
  output [31:0] io_matrixC_94_im,
  output [31:0] io_matrixC_95_re,
  output [31:0] io_matrixC_95_im,
  output [31:0] io_matrixC_96_re,
  output [31:0] io_matrixC_96_im,
  output [31:0] io_matrixC_97_re,
  output [31:0] io_matrixC_97_im,
  output [31:0] io_matrixC_98_re,
  output [31:0] io_matrixC_98_im,
  output [31:0] io_matrixC_99_re,
  output [31:0] io_matrixC_99_im,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
`endif // RANDOMIZE_REG_INIT
  wire  PE_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_1_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_1_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_1_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_1_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_1_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_1_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_1_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_1_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_1_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_1_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_1_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_1_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_2_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_2_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_2_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_2_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_2_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_2_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_2_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_2_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_2_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_2_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_2_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_2_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_3_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_3_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_3_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_3_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_3_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_3_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_3_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_3_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_3_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_3_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_3_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_3_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_4_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_4_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_4_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_4_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_4_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_4_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_4_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_4_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_4_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_4_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_4_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_4_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_5_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_5_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_5_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_5_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_5_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_5_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_5_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_5_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_5_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_5_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_5_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_5_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_6_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_6_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_6_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_6_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_6_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_6_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_6_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_6_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_6_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_6_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_6_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_6_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_7_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_7_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_7_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_7_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_7_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_7_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_7_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_7_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_7_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_7_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_7_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_7_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_8_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_8_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_8_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_8_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_8_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_8_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_8_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_8_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_8_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_8_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_8_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_8_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_9_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_9_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_9_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_9_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_9_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_9_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_9_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_9_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_9_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_9_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_9_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_9_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_10_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_10_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_10_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_10_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_10_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_10_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_10_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_10_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_10_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_10_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_10_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_10_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_11_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_11_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_11_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_11_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_11_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_11_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_11_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_11_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_11_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_11_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_11_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_11_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_12_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_12_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_12_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_12_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_12_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_12_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_12_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_12_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_12_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_12_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_12_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_12_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_13_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_13_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_13_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_13_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_13_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_13_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_13_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_13_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_13_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_13_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_13_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_13_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_14_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_14_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_14_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_14_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_14_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_14_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_14_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_14_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_14_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_14_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_14_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_14_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_15_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_15_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_15_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_15_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_15_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_15_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_15_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_15_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_15_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_15_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_15_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_15_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_16_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_16_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_16_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_16_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_16_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_16_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_16_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_16_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_16_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_16_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_16_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_16_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_17_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_17_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_17_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_17_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_17_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_17_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_17_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_17_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_17_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_17_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_17_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_17_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_18_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_18_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_18_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_18_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_18_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_18_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_18_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_18_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_18_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_18_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_18_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_18_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_19_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_19_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_19_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_19_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_19_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_19_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_19_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_19_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_19_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_19_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_19_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_19_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_20_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_20_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_20_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_20_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_20_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_20_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_20_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_20_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_20_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_20_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_20_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_20_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_21_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_21_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_21_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_21_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_21_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_21_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_21_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_21_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_21_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_21_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_21_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_21_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_22_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_22_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_22_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_22_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_22_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_22_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_22_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_22_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_22_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_22_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_22_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_22_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_23_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_23_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_23_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_23_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_23_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_23_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_23_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_23_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_23_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_23_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_23_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_23_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_24_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_24_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_24_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_24_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_24_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_24_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_24_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_24_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_24_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_24_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_24_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_24_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_25_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_25_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_25_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_25_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_25_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_25_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_25_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_25_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_25_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_25_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_25_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_25_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_26_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_26_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_26_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_26_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_26_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_26_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_26_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_26_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_26_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_26_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_26_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_26_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_27_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_27_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_27_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_27_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_27_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_27_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_27_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_27_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_27_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_27_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_27_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_27_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_28_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_28_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_28_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_28_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_28_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_28_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_28_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_28_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_28_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_28_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_28_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_28_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_29_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_29_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_29_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_29_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_29_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_29_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_29_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_29_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_29_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_29_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_29_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_29_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_30_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_30_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_30_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_30_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_30_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_30_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_30_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_30_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_30_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_30_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_30_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_30_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_31_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_31_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_31_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_31_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_31_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_31_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_31_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_31_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_31_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_31_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_31_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_31_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_32_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_32_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_32_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_32_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_32_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_32_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_32_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_32_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_32_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_32_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_32_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_32_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_33_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_33_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_33_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_33_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_33_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_33_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_33_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_33_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_33_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_33_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_33_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_33_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_34_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_34_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_34_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_34_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_34_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_34_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_34_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_34_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_34_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_34_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_34_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_34_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_35_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_35_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_35_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_35_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_35_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_35_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_35_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_35_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_35_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_35_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_35_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_35_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_36_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_36_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_36_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_36_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_36_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_36_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_36_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_36_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_36_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_36_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_36_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_36_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_37_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_37_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_37_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_37_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_37_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_37_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_37_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_37_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_37_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_37_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_37_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_37_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_38_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_38_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_38_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_38_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_38_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_38_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_38_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_38_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_38_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_38_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_38_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_38_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_39_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_39_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_39_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_39_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_39_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_39_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_39_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_39_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_39_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_39_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_39_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_39_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_40_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_40_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_40_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_40_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_40_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_40_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_40_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_40_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_40_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_40_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_40_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_40_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_41_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_41_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_41_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_41_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_41_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_41_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_41_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_41_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_41_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_41_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_41_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_41_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_42_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_42_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_42_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_42_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_42_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_42_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_42_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_42_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_42_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_42_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_42_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_42_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_43_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_43_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_43_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_43_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_43_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_43_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_43_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_43_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_43_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_43_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_43_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_43_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_44_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_44_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_44_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_44_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_44_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_44_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_44_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_44_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_44_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_44_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_44_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_44_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_45_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_45_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_45_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_45_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_45_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_45_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_45_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_45_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_45_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_45_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_45_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_45_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_46_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_46_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_46_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_46_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_46_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_46_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_46_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_46_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_46_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_46_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_46_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_46_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_47_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_47_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_47_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_47_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_47_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_47_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_47_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_47_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_47_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_47_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_47_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_47_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_48_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_48_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_48_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_48_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_48_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_48_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_48_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_48_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_48_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_48_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_48_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_48_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_49_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_49_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_49_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_49_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_49_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_49_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_49_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_49_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_49_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_49_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_49_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_49_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_50_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_50_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_50_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_50_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_50_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_50_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_50_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_50_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_50_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_50_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_50_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_50_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_51_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_51_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_51_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_51_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_51_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_51_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_51_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_51_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_51_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_51_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_51_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_51_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_52_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_52_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_52_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_52_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_52_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_52_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_52_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_52_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_52_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_52_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_52_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_52_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_53_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_53_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_53_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_53_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_53_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_53_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_53_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_53_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_53_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_53_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_53_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_53_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_54_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_54_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_54_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_54_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_54_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_54_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_54_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_54_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_54_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_54_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_54_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_54_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_55_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_55_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_55_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_55_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_55_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_55_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_55_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_55_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_55_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_55_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_55_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_55_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_56_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_56_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_56_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_56_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_56_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_56_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_56_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_56_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_56_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_56_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_56_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_56_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_57_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_57_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_57_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_57_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_57_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_57_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_57_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_57_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_57_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_57_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_57_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_57_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_58_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_58_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_58_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_58_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_58_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_58_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_58_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_58_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_58_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_58_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_58_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_58_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_59_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_59_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_59_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_59_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_59_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_59_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_59_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_59_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_59_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_59_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_59_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_59_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_60_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_60_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_60_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_60_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_60_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_60_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_60_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_60_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_60_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_60_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_60_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_60_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_61_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_61_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_61_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_61_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_61_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_61_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_61_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_61_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_61_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_61_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_61_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_61_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_62_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_62_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_62_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_62_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_62_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_62_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_62_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_62_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_62_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_62_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_62_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_62_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_63_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_63_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_63_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_63_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_63_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_63_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_63_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_63_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_63_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_63_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_63_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_63_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_64_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_64_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_64_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_64_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_64_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_64_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_64_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_64_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_64_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_64_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_64_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_64_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_65_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_65_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_65_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_65_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_65_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_65_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_65_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_65_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_65_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_65_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_65_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_65_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_66_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_66_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_66_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_66_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_66_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_66_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_66_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_66_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_66_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_66_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_66_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_66_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_67_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_67_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_67_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_67_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_67_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_67_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_67_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_67_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_67_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_67_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_67_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_67_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_68_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_68_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_68_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_68_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_68_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_68_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_68_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_68_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_68_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_68_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_68_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_68_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_69_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_69_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_69_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_69_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_69_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_69_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_69_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_69_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_69_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_69_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_69_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_69_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_70_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_70_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_70_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_70_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_70_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_70_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_70_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_70_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_70_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_70_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_70_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_70_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_71_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_71_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_71_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_71_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_71_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_71_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_71_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_71_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_71_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_71_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_71_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_71_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_72_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_72_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_72_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_72_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_72_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_72_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_72_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_72_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_72_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_72_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_72_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_72_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_73_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_73_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_73_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_73_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_73_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_73_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_73_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_73_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_73_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_73_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_73_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_73_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_74_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_74_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_74_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_74_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_74_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_74_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_74_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_74_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_74_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_74_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_74_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_74_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_75_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_75_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_75_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_75_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_75_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_75_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_75_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_75_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_75_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_75_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_75_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_75_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_76_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_76_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_76_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_76_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_76_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_76_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_76_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_76_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_76_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_76_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_76_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_76_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_77_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_77_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_77_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_77_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_77_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_77_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_77_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_77_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_77_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_77_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_77_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_77_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_78_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_78_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_78_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_78_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_78_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_78_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_78_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_78_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_78_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_78_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_78_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_78_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_79_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_79_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_79_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_79_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_79_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_79_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_79_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_79_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_79_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_79_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_79_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_79_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_80_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_80_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_80_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_80_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_80_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_80_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_80_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_80_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_80_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_80_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_80_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_80_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_81_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_81_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_81_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_81_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_81_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_81_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_81_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_81_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_81_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_81_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_81_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_81_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_82_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_82_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_82_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_82_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_82_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_82_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_82_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_82_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_82_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_82_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_82_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_82_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_83_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_83_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_83_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_83_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_83_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_83_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_83_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_83_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_83_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_83_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_83_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_83_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_84_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_84_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_84_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_84_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_84_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_84_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_84_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_84_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_84_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_84_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_84_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_84_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_85_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_85_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_85_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_85_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_85_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_85_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_85_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_85_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_85_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_85_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_85_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_85_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_86_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_86_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_86_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_86_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_86_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_86_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_86_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_86_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_86_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_86_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_86_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_86_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_87_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_87_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_87_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_87_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_87_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_87_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_87_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_87_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_87_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_87_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_87_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_87_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_88_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_88_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_88_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_88_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_88_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_88_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_88_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_88_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_88_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_88_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_88_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_88_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_89_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_89_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_89_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_89_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_89_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_89_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_89_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_89_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_89_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_89_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_89_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_89_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_90_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_90_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_90_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_90_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_90_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_90_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_90_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_90_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_90_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_90_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_90_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_90_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_91_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_91_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_91_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_91_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_91_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_91_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_91_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_91_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_91_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_91_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_91_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_91_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_92_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_92_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_92_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_92_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_92_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_92_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_92_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_92_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_92_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_92_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_92_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_92_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_93_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_93_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_93_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_93_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_93_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_93_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_93_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_93_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_93_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_93_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_93_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_93_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_94_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_94_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_94_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_94_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_94_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_94_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_94_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_94_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_94_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_94_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_94_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_94_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_95_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_95_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_95_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_95_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_95_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_95_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_95_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_95_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_95_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_95_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_95_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_95_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_96_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_96_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_96_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_96_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_96_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_96_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_96_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_96_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_96_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_96_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_96_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_96_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_97_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_97_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_97_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_97_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_97_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_97_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_97_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_97_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_97_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_97_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_97_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_97_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_98_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_98_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_98_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_98_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_98_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_98_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_98_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_98_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_98_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_98_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_98_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_98_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_99_clock; // @[Matrix_Mul_V1.scala 86:35]
  wire  PE_99_io_reset; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_99_io_in_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_99_io_in_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_99_io_in_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_99_io_in_y_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_99_io_out_pe_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_99_io_out_pe_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_99_io_out_x_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_99_io_out_x_im; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_99_io_out_y_re; // @[Matrix_Mul_V1.scala 86:35]
  wire [31:0] PE_99_io_out_y_im; // @[Matrix_Mul_V1.scala 86:35]
  reg [31:0] regsA_0_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_0_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_1_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_1_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_2_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_2_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_3_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_3_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_4_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_4_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_5_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_5_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_6_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_6_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_7_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_7_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_8_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_8_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_9_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_9_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_10_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_10_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_11_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_11_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_12_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_12_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_13_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_13_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_14_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_14_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_15_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_15_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_16_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_16_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_17_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_17_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_18_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_18_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_19_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_19_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_20_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_20_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_21_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_21_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_22_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_22_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_23_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_23_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_24_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_24_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_25_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_25_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_26_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_26_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_27_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_27_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_28_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_28_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_29_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_29_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_30_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_30_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_31_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_31_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_32_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_32_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_33_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_33_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_34_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_34_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_35_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_35_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_36_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_36_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_37_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_37_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_38_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_38_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_39_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_39_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_40_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_40_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_41_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_41_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_42_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_42_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_43_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_43_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_44_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_44_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_45_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_45_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_46_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_46_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_47_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_47_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_48_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_48_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_49_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_49_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_50_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_50_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_51_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_51_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_52_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_52_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_53_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_53_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_54_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_54_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_55_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_55_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_56_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_56_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_57_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_57_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_58_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_58_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_59_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_59_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_60_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_60_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_61_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_61_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_62_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_62_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_63_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_63_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_64_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_64_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_65_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_65_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_66_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_66_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_67_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_67_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_68_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_68_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_69_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_69_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_70_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_70_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_71_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_71_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_72_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_72_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_73_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_73_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_74_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_74_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_75_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_75_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_76_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_76_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_77_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_77_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_78_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_78_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_79_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_79_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_80_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_80_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_81_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_81_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_82_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_82_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_83_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_83_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_84_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_84_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_85_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_85_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_86_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_86_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_87_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_87_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_88_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_88_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_89_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_89_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_90_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_90_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_91_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_91_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_92_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_92_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_93_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_93_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_94_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_94_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_95_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_95_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_96_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_96_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_97_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_97_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_98_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_98_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_99_re; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsA_99_im; // @[Matrix_Mul_V1.scala 82:32]
  reg [31:0] regsB_0_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_0_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_1_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_1_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_2_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_2_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_3_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_3_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_4_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_4_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_5_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_5_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_6_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_6_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_7_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_7_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_8_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_8_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_9_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_9_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_10_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_10_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_11_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_11_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_12_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_12_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_13_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_13_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_14_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_14_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_15_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_15_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_16_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_16_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_17_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_17_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_18_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_18_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_19_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_19_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_20_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_20_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_21_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_21_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_22_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_22_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_23_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_23_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_24_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_24_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_25_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_25_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_26_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_26_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_27_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_27_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_28_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_28_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_29_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_29_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_30_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_30_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_31_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_31_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_32_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_32_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_33_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_33_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_34_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_34_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_35_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_35_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_36_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_36_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_37_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_37_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_38_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_38_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_39_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_39_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_40_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_40_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_41_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_41_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_42_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_42_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_43_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_43_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_44_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_44_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_45_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_45_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_46_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_46_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_47_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_47_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_48_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_48_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_49_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_49_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_50_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_50_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_51_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_51_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_52_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_52_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_53_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_53_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_54_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_54_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_55_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_55_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_56_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_56_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_57_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_57_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_58_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_58_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_59_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_59_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_60_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_60_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_61_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_61_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_62_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_62_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_63_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_63_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_64_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_64_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_65_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_65_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_66_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_66_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_67_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_67_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_68_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_68_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_69_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_69_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_70_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_70_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_71_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_71_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_72_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_72_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_73_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_73_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_74_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_74_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_75_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_75_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_76_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_76_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_77_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_77_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_78_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_78_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_79_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_79_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_80_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_80_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_81_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_81_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_82_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_82_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_83_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_83_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_84_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_84_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_85_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_85_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_86_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_86_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_87_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_87_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_88_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_88_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_89_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_89_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_90_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_90_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_91_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_91_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_92_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_92_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_93_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_93_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_94_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_94_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_95_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_95_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_96_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_96_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_97_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_97_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_98_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_98_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_99_re; // @[Matrix_Mul_V1.scala 83:32]
  reg [31:0] regsB_99_im; // @[Matrix_Mul_V1.scala 83:32]
  reg [5:0] input_point; // @[Matrix_Mul_V1.scala 84:30]
  wire [5:0] _input_point_T_1 = input_point + 6'h1; // @[Matrix_Mul_V1.scala 116:32]
  wire  _T = input_point < 6'h13; // @[Matrix_Mul_V1.scala 145:20]
  wire [5:0] _T_1 = 1'h0 * 5'h13; // @[Matrix_Mul_V1.scala 148:44]
  wire [5:0] _T_3 = _T_1 + input_point; // @[Matrix_Mul_V1.scala 148:60]
  wire [31:0] _GEN_805 = 6'h1 == _T_3 ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_806 = 6'h2 == _T_3 ? $signed(regsA_2_im) : $signed(_GEN_805); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_807 = 6'h3 == _T_3 ? $signed(regsA_3_im) : $signed(_GEN_806); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_808 = 6'h4 == _T_3 ? $signed(regsA_4_im) : $signed(_GEN_807); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_809 = 6'h5 == _T_3 ? $signed(regsA_5_im) : $signed(_GEN_808); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_810 = 6'h6 == _T_3 ? $signed(regsA_6_im) : $signed(_GEN_809); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_811 = 6'h7 == _T_3 ? $signed(regsA_7_im) : $signed(_GEN_810); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_812 = 6'h8 == _T_3 ? $signed(regsA_8_im) : $signed(_GEN_811); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_813 = 6'h9 == _T_3 ? $signed(regsA_9_im) : $signed(_GEN_812); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_814 = 6'ha == _T_3 ? $signed(32'sh0) : $signed(_GEN_813); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_815 = 6'hb == _T_3 ? $signed(32'sh0) : $signed(_GEN_814); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_816 = 6'hc == _T_3 ? $signed(32'sh0) : $signed(_GEN_815); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_817 = 6'hd == _T_3 ? $signed(32'sh0) : $signed(_GEN_816); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_818 = 6'he == _T_3 ? $signed(32'sh0) : $signed(_GEN_817); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_819 = 6'hf == _T_3 ? $signed(32'sh0) : $signed(_GEN_818); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_820 = 6'h10 == _T_3 ? $signed(32'sh0) : $signed(_GEN_819); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_821 = 6'h11 == _T_3 ? $signed(32'sh0) : $signed(_GEN_820); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_822 = 6'h12 == _T_3 ? $signed(32'sh0) : $signed(_GEN_821); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_823 = 6'h13 == _T_3 ? $signed(32'sh0) : $signed(_GEN_822); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_824 = 6'h14 == _T_3 ? $signed(regsA_10_im) : $signed(_GEN_823); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_825 = 6'h15 == _T_3 ? $signed(regsA_11_im) : $signed(_GEN_824); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_826 = 6'h16 == _T_3 ? $signed(regsA_12_im) : $signed(_GEN_825); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_827 = 6'h17 == _T_3 ? $signed(regsA_13_im) : $signed(_GEN_826); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_828 = 6'h18 == _T_3 ? $signed(regsA_14_im) : $signed(_GEN_827); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_829 = 6'h19 == _T_3 ? $signed(regsA_15_im) : $signed(_GEN_828); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_830 = 6'h1a == _T_3 ? $signed(regsA_16_im) : $signed(_GEN_829); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_831 = 6'h1b == _T_3 ? $signed(regsA_17_im) : $signed(_GEN_830); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_832 = 6'h1c == _T_3 ? $signed(regsA_18_im) : $signed(_GEN_831); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_833 = 6'h1d == _T_3 ? $signed(regsA_19_im) : $signed(_GEN_832); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_834 = 6'h1e == _T_3 ? $signed(32'sh0) : $signed(_GEN_833); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_835 = 6'h1f == _T_3 ? $signed(32'sh0) : $signed(_GEN_834); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_836 = 6'h20 == _T_3 ? $signed(32'sh0) : $signed(_GEN_835); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_837 = 6'h21 == _T_3 ? $signed(32'sh0) : $signed(_GEN_836); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_838 = 6'h22 == _T_3 ? $signed(32'sh0) : $signed(_GEN_837); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_839 = 6'h23 == _T_3 ? $signed(32'sh0) : $signed(_GEN_838); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_840 = 6'h24 == _T_3 ? $signed(32'sh0) : $signed(_GEN_839); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_841 = 6'h25 == _T_3 ? $signed(32'sh0) : $signed(_GEN_840); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_842 = 6'h26 == _T_3 ? $signed(32'sh0) : $signed(_GEN_841); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_843 = 6'h27 == _T_3 ? $signed(32'sh0) : $signed(_GEN_842); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_844 = 6'h28 == _T_3 ? $signed(regsA_20_im) : $signed(_GEN_843); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_845 = 6'h29 == _T_3 ? $signed(regsA_21_im) : $signed(_GEN_844); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_846 = 6'h2a == _T_3 ? $signed(regsA_22_im) : $signed(_GEN_845); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_847 = 6'h2b == _T_3 ? $signed(regsA_23_im) : $signed(_GEN_846); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_848 = 6'h2c == _T_3 ? $signed(regsA_24_im) : $signed(_GEN_847); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_849 = 6'h2d == _T_3 ? $signed(regsA_25_im) : $signed(_GEN_848); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_850 = 6'h2e == _T_3 ? $signed(regsA_26_im) : $signed(_GEN_849); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_851 = 6'h2f == _T_3 ? $signed(regsA_27_im) : $signed(_GEN_850); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_852 = 6'h30 == _T_3 ? $signed(regsA_28_im) : $signed(_GEN_851); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_853 = 6'h31 == _T_3 ? $signed(regsA_29_im) : $signed(_GEN_852); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_854 = 6'h32 == _T_3 ? $signed(32'sh0) : $signed(_GEN_853); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_855 = 6'h33 == _T_3 ? $signed(32'sh0) : $signed(_GEN_854); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_856 = 6'h34 == _T_3 ? $signed(32'sh0) : $signed(_GEN_855); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_857 = 6'h35 == _T_3 ? $signed(32'sh0) : $signed(_GEN_856); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_858 = 6'h36 == _T_3 ? $signed(32'sh0) : $signed(_GEN_857); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_859 = 6'h37 == _T_3 ? $signed(32'sh0) : $signed(_GEN_858); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_860 = 6'h38 == _T_3 ? $signed(32'sh0) : $signed(_GEN_859); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_861 = 6'h39 == _T_3 ? $signed(32'sh0) : $signed(_GEN_860); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_862 = 6'h3a == _T_3 ? $signed(32'sh0) : $signed(_GEN_861); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_863 = 6'h3b == _T_3 ? $signed(32'sh0) : $signed(_GEN_862); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_864 = 6'h3c == _T_3 ? $signed(regsA_30_im) : $signed(_GEN_863); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_865 = 6'h3d == _T_3 ? $signed(regsA_31_im) : $signed(_GEN_864); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_866 = 6'h3e == _T_3 ? $signed(regsA_32_im) : $signed(_GEN_865); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_867 = 6'h3f == _T_3 ? $signed(regsA_33_im) : $signed(_GEN_866); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [6:0] _GEN_8445 = {{1'd0}, _T_3}; // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_868 = 7'h40 == _GEN_8445 ? $signed(regsA_34_im) : $signed(_GEN_867); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_869 = 7'h41 == _GEN_8445 ? $signed(regsA_35_im) : $signed(_GEN_868); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_870 = 7'h42 == _GEN_8445 ? $signed(regsA_36_im) : $signed(_GEN_869); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_871 = 7'h43 == _GEN_8445 ? $signed(regsA_37_im) : $signed(_GEN_870); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_872 = 7'h44 == _GEN_8445 ? $signed(regsA_38_im) : $signed(_GEN_871); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_873 = 7'h45 == _GEN_8445 ? $signed(regsA_39_im) : $signed(_GEN_872); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_874 = 7'h46 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_873); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_875 = 7'h47 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_874); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_876 = 7'h48 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_875); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_877 = 7'h49 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_876); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_878 = 7'h4a == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_877); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_879 = 7'h4b == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_878); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_880 = 7'h4c == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_879); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_881 = 7'h4d == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_880); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_882 = 7'h4e == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_881); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_883 = 7'h4f == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_882); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_884 = 7'h50 == _GEN_8445 ? $signed(regsA_40_im) : $signed(_GEN_883); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_885 = 7'h51 == _GEN_8445 ? $signed(regsA_41_im) : $signed(_GEN_884); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_886 = 7'h52 == _GEN_8445 ? $signed(regsA_42_im) : $signed(_GEN_885); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_887 = 7'h53 == _GEN_8445 ? $signed(regsA_43_im) : $signed(_GEN_886); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_888 = 7'h54 == _GEN_8445 ? $signed(regsA_44_im) : $signed(_GEN_887); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_889 = 7'h55 == _GEN_8445 ? $signed(regsA_45_im) : $signed(_GEN_888); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_890 = 7'h56 == _GEN_8445 ? $signed(regsA_46_im) : $signed(_GEN_889); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_891 = 7'h57 == _GEN_8445 ? $signed(regsA_47_im) : $signed(_GEN_890); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_892 = 7'h58 == _GEN_8445 ? $signed(regsA_48_im) : $signed(_GEN_891); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_893 = 7'h59 == _GEN_8445 ? $signed(regsA_49_im) : $signed(_GEN_892); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_894 = 7'h5a == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_893); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_895 = 7'h5b == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_894); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_896 = 7'h5c == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_895); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_897 = 7'h5d == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_896); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_898 = 7'h5e == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_897); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_899 = 7'h5f == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_898); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_900 = 7'h60 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_899); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_901 = 7'h61 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_900); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_902 = 7'h62 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_901); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_903 = 7'h63 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_902); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_904 = 7'h64 == _GEN_8445 ? $signed(regsA_50_im) : $signed(_GEN_903); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_905 = 7'h65 == _GEN_8445 ? $signed(regsA_51_im) : $signed(_GEN_904); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_906 = 7'h66 == _GEN_8445 ? $signed(regsA_52_im) : $signed(_GEN_905); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_907 = 7'h67 == _GEN_8445 ? $signed(regsA_53_im) : $signed(_GEN_906); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_908 = 7'h68 == _GEN_8445 ? $signed(regsA_54_im) : $signed(_GEN_907); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_909 = 7'h69 == _GEN_8445 ? $signed(regsA_55_im) : $signed(_GEN_908); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_910 = 7'h6a == _GEN_8445 ? $signed(regsA_56_im) : $signed(_GEN_909); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_911 = 7'h6b == _GEN_8445 ? $signed(regsA_57_im) : $signed(_GEN_910); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_912 = 7'h6c == _GEN_8445 ? $signed(regsA_58_im) : $signed(_GEN_911); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_913 = 7'h6d == _GEN_8445 ? $signed(regsA_59_im) : $signed(_GEN_912); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_914 = 7'h6e == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_913); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_915 = 7'h6f == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_914); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_916 = 7'h70 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_915); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_917 = 7'h71 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_916); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_918 = 7'h72 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_917); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_919 = 7'h73 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_918); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_920 = 7'h74 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_919); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_921 = 7'h75 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_920); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_922 = 7'h76 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_921); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_923 = 7'h77 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_922); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_924 = 7'h78 == _GEN_8445 ? $signed(regsA_60_im) : $signed(_GEN_923); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_925 = 7'h79 == _GEN_8445 ? $signed(regsA_61_im) : $signed(_GEN_924); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_926 = 7'h7a == _GEN_8445 ? $signed(regsA_62_im) : $signed(_GEN_925); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_927 = 7'h7b == _GEN_8445 ? $signed(regsA_63_im) : $signed(_GEN_926); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_928 = 7'h7c == _GEN_8445 ? $signed(regsA_64_im) : $signed(_GEN_927); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_929 = 7'h7d == _GEN_8445 ? $signed(regsA_65_im) : $signed(_GEN_928); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_930 = 7'h7e == _GEN_8445 ? $signed(regsA_66_im) : $signed(_GEN_929); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_931 = 7'h7f == _GEN_8445 ? $signed(regsA_67_im) : $signed(_GEN_930); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [7:0] _GEN_8509 = {{2'd0}, _T_3}; // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_932 = 8'h80 == _GEN_8509 ? $signed(regsA_68_im) : $signed(_GEN_931); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_933 = 8'h81 == _GEN_8509 ? $signed(regsA_69_im) : $signed(_GEN_932); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_934 = 8'h82 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_933); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_935 = 8'h83 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_934); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_936 = 8'h84 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_935); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_937 = 8'h85 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_936); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_938 = 8'h86 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_937); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_939 = 8'h87 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_938); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_940 = 8'h88 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_939); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_941 = 8'h89 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_940); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_942 = 8'h8a == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_941); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_943 = 8'h8b == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_942); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_944 = 8'h8c == _GEN_8509 ? $signed(regsA_70_im) : $signed(_GEN_943); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_945 = 8'h8d == _GEN_8509 ? $signed(regsA_71_im) : $signed(_GEN_944); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_946 = 8'h8e == _GEN_8509 ? $signed(regsA_72_im) : $signed(_GEN_945); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_947 = 8'h8f == _GEN_8509 ? $signed(regsA_73_im) : $signed(_GEN_946); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_948 = 8'h90 == _GEN_8509 ? $signed(regsA_74_im) : $signed(_GEN_947); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_949 = 8'h91 == _GEN_8509 ? $signed(regsA_75_im) : $signed(_GEN_948); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_950 = 8'h92 == _GEN_8509 ? $signed(regsA_76_im) : $signed(_GEN_949); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_951 = 8'h93 == _GEN_8509 ? $signed(regsA_77_im) : $signed(_GEN_950); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_952 = 8'h94 == _GEN_8509 ? $signed(regsA_78_im) : $signed(_GEN_951); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_953 = 8'h95 == _GEN_8509 ? $signed(regsA_79_im) : $signed(_GEN_952); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_954 = 8'h96 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_953); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_955 = 8'h97 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_954); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_956 = 8'h98 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_955); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_957 = 8'h99 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_956); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_958 = 8'h9a == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_957); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_959 = 8'h9b == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_958); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_960 = 8'h9c == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_959); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_961 = 8'h9d == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_960); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_962 = 8'h9e == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_961); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_963 = 8'h9f == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_962); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_964 = 8'ha0 == _GEN_8509 ? $signed(regsA_80_im) : $signed(_GEN_963); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_965 = 8'ha1 == _GEN_8509 ? $signed(regsA_81_im) : $signed(_GEN_964); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_966 = 8'ha2 == _GEN_8509 ? $signed(regsA_82_im) : $signed(_GEN_965); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_967 = 8'ha3 == _GEN_8509 ? $signed(regsA_83_im) : $signed(_GEN_966); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_968 = 8'ha4 == _GEN_8509 ? $signed(regsA_84_im) : $signed(_GEN_967); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_969 = 8'ha5 == _GEN_8509 ? $signed(regsA_85_im) : $signed(_GEN_968); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_970 = 8'ha6 == _GEN_8509 ? $signed(regsA_86_im) : $signed(_GEN_969); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_971 = 8'ha7 == _GEN_8509 ? $signed(regsA_87_im) : $signed(_GEN_970); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_972 = 8'ha8 == _GEN_8509 ? $signed(regsA_88_im) : $signed(_GEN_971); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_973 = 8'ha9 == _GEN_8509 ? $signed(regsA_89_im) : $signed(_GEN_972); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_974 = 8'haa == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_973); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_975 = 8'hab == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_974); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_976 = 8'hac == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_975); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_977 = 8'had == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_976); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_978 = 8'hae == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_977); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_979 = 8'haf == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_978); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_980 = 8'hb0 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_979); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_981 = 8'hb1 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_980); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_982 = 8'hb2 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_981); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_983 = 8'hb3 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_982); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_984 = 8'hb4 == _GEN_8509 ? $signed(regsA_90_im) : $signed(_GEN_983); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_985 = 8'hb5 == _GEN_8509 ? $signed(regsA_91_im) : $signed(_GEN_984); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_986 = 8'hb6 == _GEN_8509 ? $signed(regsA_92_im) : $signed(_GEN_985); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_987 = 8'hb7 == _GEN_8509 ? $signed(regsA_93_im) : $signed(_GEN_986); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_988 = 8'hb8 == _GEN_8509 ? $signed(regsA_94_im) : $signed(_GEN_987); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_989 = 8'hb9 == _GEN_8509 ? $signed(regsA_95_im) : $signed(_GEN_988); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_990 = 8'hba == _GEN_8509 ? $signed(regsA_96_im) : $signed(_GEN_989); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_991 = 8'hbb == _GEN_8509 ? $signed(regsA_97_im) : $signed(_GEN_990); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_992 = 8'hbc == _GEN_8509 ? $signed(regsA_98_im) : $signed(_GEN_991); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_993 = 8'hbd == _GEN_8509 ? $signed(regsA_99_im) : $signed(_GEN_992); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_995 = 6'h1 == _T_3 ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_996 = 6'h2 == _T_3 ? $signed(regsA_2_re) : $signed(_GEN_995); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_997 = 6'h3 == _T_3 ? $signed(regsA_3_re) : $signed(_GEN_996); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_998 = 6'h4 == _T_3 ? $signed(regsA_4_re) : $signed(_GEN_997); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_999 = 6'h5 == _T_3 ? $signed(regsA_5_re) : $signed(_GEN_998); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1000 = 6'h6 == _T_3 ? $signed(regsA_6_re) : $signed(_GEN_999); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1001 = 6'h7 == _T_3 ? $signed(regsA_7_re) : $signed(_GEN_1000); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1002 = 6'h8 == _T_3 ? $signed(regsA_8_re) : $signed(_GEN_1001); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1003 = 6'h9 == _T_3 ? $signed(regsA_9_re) : $signed(_GEN_1002); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1004 = 6'ha == _T_3 ? $signed(32'sh0) : $signed(_GEN_1003); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1005 = 6'hb == _T_3 ? $signed(32'sh0) : $signed(_GEN_1004); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1006 = 6'hc == _T_3 ? $signed(32'sh0) : $signed(_GEN_1005); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1007 = 6'hd == _T_3 ? $signed(32'sh0) : $signed(_GEN_1006); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1008 = 6'he == _T_3 ? $signed(32'sh0) : $signed(_GEN_1007); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1009 = 6'hf == _T_3 ? $signed(32'sh0) : $signed(_GEN_1008); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1010 = 6'h10 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1009); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1011 = 6'h11 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1010); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1012 = 6'h12 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1011); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1013 = 6'h13 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1012); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1014 = 6'h14 == _T_3 ? $signed(regsA_10_re) : $signed(_GEN_1013); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1015 = 6'h15 == _T_3 ? $signed(regsA_11_re) : $signed(_GEN_1014); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1016 = 6'h16 == _T_3 ? $signed(regsA_12_re) : $signed(_GEN_1015); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1017 = 6'h17 == _T_3 ? $signed(regsA_13_re) : $signed(_GEN_1016); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1018 = 6'h18 == _T_3 ? $signed(regsA_14_re) : $signed(_GEN_1017); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1019 = 6'h19 == _T_3 ? $signed(regsA_15_re) : $signed(_GEN_1018); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1020 = 6'h1a == _T_3 ? $signed(regsA_16_re) : $signed(_GEN_1019); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1021 = 6'h1b == _T_3 ? $signed(regsA_17_re) : $signed(_GEN_1020); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1022 = 6'h1c == _T_3 ? $signed(regsA_18_re) : $signed(_GEN_1021); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1023 = 6'h1d == _T_3 ? $signed(regsA_19_re) : $signed(_GEN_1022); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1024 = 6'h1e == _T_3 ? $signed(32'sh0) : $signed(_GEN_1023); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1025 = 6'h1f == _T_3 ? $signed(32'sh0) : $signed(_GEN_1024); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1026 = 6'h20 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1025); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1027 = 6'h21 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1026); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1028 = 6'h22 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1027); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1029 = 6'h23 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1028); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1030 = 6'h24 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1029); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1031 = 6'h25 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1030); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1032 = 6'h26 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1031); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1033 = 6'h27 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1032); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1034 = 6'h28 == _T_3 ? $signed(regsA_20_re) : $signed(_GEN_1033); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1035 = 6'h29 == _T_3 ? $signed(regsA_21_re) : $signed(_GEN_1034); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1036 = 6'h2a == _T_3 ? $signed(regsA_22_re) : $signed(_GEN_1035); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1037 = 6'h2b == _T_3 ? $signed(regsA_23_re) : $signed(_GEN_1036); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1038 = 6'h2c == _T_3 ? $signed(regsA_24_re) : $signed(_GEN_1037); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1039 = 6'h2d == _T_3 ? $signed(regsA_25_re) : $signed(_GEN_1038); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1040 = 6'h2e == _T_3 ? $signed(regsA_26_re) : $signed(_GEN_1039); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1041 = 6'h2f == _T_3 ? $signed(regsA_27_re) : $signed(_GEN_1040); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1042 = 6'h30 == _T_3 ? $signed(regsA_28_re) : $signed(_GEN_1041); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1043 = 6'h31 == _T_3 ? $signed(regsA_29_re) : $signed(_GEN_1042); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1044 = 6'h32 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1043); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1045 = 6'h33 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1044); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1046 = 6'h34 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1045); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1047 = 6'h35 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1046); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1048 = 6'h36 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1047); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1049 = 6'h37 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1048); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1050 = 6'h38 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1049); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1051 = 6'h39 == _T_3 ? $signed(32'sh0) : $signed(_GEN_1050); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1052 = 6'h3a == _T_3 ? $signed(32'sh0) : $signed(_GEN_1051); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1053 = 6'h3b == _T_3 ? $signed(32'sh0) : $signed(_GEN_1052); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1054 = 6'h3c == _T_3 ? $signed(regsA_30_re) : $signed(_GEN_1053); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1055 = 6'h3d == _T_3 ? $signed(regsA_31_re) : $signed(_GEN_1054); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1056 = 6'h3e == _T_3 ? $signed(regsA_32_re) : $signed(_GEN_1055); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1057 = 6'h3f == _T_3 ? $signed(regsA_33_re) : $signed(_GEN_1056); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1058 = 7'h40 == _GEN_8445 ? $signed(regsA_34_re) : $signed(_GEN_1057); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1059 = 7'h41 == _GEN_8445 ? $signed(regsA_35_re) : $signed(_GEN_1058); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1060 = 7'h42 == _GEN_8445 ? $signed(regsA_36_re) : $signed(_GEN_1059); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1061 = 7'h43 == _GEN_8445 ? $signed(regsA_37_re) : $signed(_GEN_1060); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1062 = 7'h44 == _GEN_8445 ? $signed(regsA_38_re) : $signed(_GEN_1061); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1063 = 7'h45 == _GEN_8445 ? $signed(regsA_39_re) : $signed(_GEN_1062); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1064 = 7'h46 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1063); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1065 = 7'h47 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1064); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1066 = 7'h48 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1065); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1067 = 7'h49 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1066); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1068 = 7'h4a == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1067); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1069 = 7'h4b == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1068); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1070 = 7'h4c == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1069); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1071 = 7'h4d == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1070); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1072 = 7'h4e == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1071); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1073 = 7'h4f == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1072); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1074 = 7'h50 == _GEN_8445 ? $signed(regsA_40_re) : $signed(_GEN_1073); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1075 = 7'h51 == _GEN_8445 ? $signed(regsA_41_re) : $signed(_GEN_1074); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1076 = 7'h52 == _GEN_8445 ? $signed(regsA_42_re) : $signed(_GEN_1075); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1077 = 7'h53 == _GEN_8445 ? $signed(regsA_43_re) : $signed(_GEN_1076); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1078 = 7'h54 == _GEN_8445 ? $signed(regsA_44_re) : $signed(_GEN_1077); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1079 = 7'h55 == _GEN_8445 ? $signed(regsA_45_re) : $signed(_GEN_1078); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1080 = 7'h56 == _GEN_8445 ? $signed(regsA_46_re) : $signed(_GEN_1079); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1081 = 7'h57 == _GEN_8445 ? $signed(regsA_47_re) : $signed(_GEN_1080); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1082 = 7'h58 == _GEN_8445 ? $signed(regsA_48_re) : $signed(_GEN_1081); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1083 = 7'h59 == _GEN_8445 ? $signed(regsA_49_re) : $signed(_GEN_1082); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1084 = 7'h5a == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1083); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1085 = 7'h5b == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1084); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1086 = 7'h5c == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1085); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1087 = 7'h5d == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1086); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1088 = 7'h5e == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1087); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1089 = 7'h5f == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1088); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1090 = 7'h60 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1089); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1091 = 7'h61 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1090); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1092 = 7'h62 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1091); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1093 = 7'h63 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1092); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1094 = 7'h64 == _GEN_8445 ? $signed(regsA_50_re) : $signed(_GEN_1093); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1095 = 7'h65 == _GEN_8445 ? $signed(regsA_51_re) : $signed(_GEN_1094); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1096 = 7'h66 == _GEN_8445 ? $signed(regsA_52_re) : $signed(_GEN_1095); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1097 = 7'h67 == _GEN_8445 ? $signed(regsA_53_re) : $signed(_GEN_1096); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1098 = 7'h68 == _GEN_8445 ? $signed(regsA_54_re) : $signed(_GEN_1097); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1099 = 7'h69 == _GEN_8445 ? $signed(regsA_55_re) : $signed(_GEN_1098); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1100 = 7'h6a == _GEN_8445 ? $signed(regsA_56_re) : $signed(_GEN_1099); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1101 = 7'h6b == _GEN_8445 ? $signed(regsA_57_re) : $signed(_GEN_1100); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1102 = 7'h6c == _GEN_8445 ? $signed(regsA_58_re) : $signed(_GEN_1101); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1103 = 7'h6d == _GEN_8445 ? $signed(regsA_59_re) : $signed(_GEN_1102); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1104 = 7'h6e == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1103); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1105 = 7'h6f == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1104); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1106 = 7'h70 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1105); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1107 = 7'h71 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1106); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1108 = 7'h72 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1107); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1109 = 7'h73 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1108); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1110 = 7'h74 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1109); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1111 = 7'h75 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1110); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1112 = 7'h76 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1111); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1113 = 7'h77 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_1112); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1114 = 7'h78 == _GEN_8445 ? $signed(regsA_60_re) : $signed(_GEN_1113); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1115 = 7'h79 == _GEN_8445 ? $signed(regsA_61_re) : $signed(_GEN_1114); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1116 = 7'h7a == _GEN_8445 ? $signed(regsA_62_re) : $signed(_GEN_1115); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1117 = 7'h7b == _GEN_8445 ? $signed(regsA_63_re) : $signed(_GEN_1116); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1118 = 7'h7c == _GEN_8445 ? $signed(regsA_64_re) : $signed(_GEN_1117); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1119 = 7'h7d == _GEN_8445 ? $signed(regsA_65_re) : $signed(_GEN_1118); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1120 = 7'h7e == _GEN_8445 ? $signed(regsA_66_re) : $signed(_GEN_1119); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1121 = 7'h7f == _GEN_8445 ? $signed(regsA_67_re) : $signed(_GEN_1120); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1122 = 8'h80 == _GEN_8509 ? $signed(regsA_68_re) : $signed(_GEN_1121); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1123 = 8'h81 == _GEN_8509 ? $signed(regsA_69_re) : $signed(_GEN_1122); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1124 = 8'h82 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1123); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1125 = 8'h83 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1124); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1126 = 8'h84 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1125); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1127 = 8'h85 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1126); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1128 = 8'h86 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1127); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1129 = 8'h87 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1128); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1130 = 8'h88 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1129); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1131 = 8'h89 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1130); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1132 = 8'h8a == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1131); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1133 = 8'h8b == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1132); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1134 = 8'h8c == _GEN_8509 ? $signed(regsA_70_re) : $signed(_GEN_1133); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1135 = 8'h8d == _GEN_8509 ? $signed(regsA_71_re) : $signed(_GEN_1134); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1136 = 8'h8e == _GEN_8509 ? $signed(regsA_72_re) : $signed(_GEN_1135); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1137 = 8'h8f == _GEN_8509 ? $signed(regsA_73_re) : $signed(_GEN_1136); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1138 = 8'h90 == _GEN_8509 ? $signed(regsA_74_re) : $signed(_GEN_1137); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1139 = 8'h91 == _GEN_8509 ? $signed(regsA_75_re) : $signed(_GEN_1138); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1140 = 8'h92 == _GEN_8509 ? $signed(regsA_76_re) : $signed(_GEN_1139); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1141 = 8'h93 == _GEN_8509 ? $signed(regsA_77_re) : $signed(_GEN_1140); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1142 = 8'h94 == _GEN_8509 ? $signed(regsA_78_re) : $signed(_GEN_1141); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1143 = 8'h95 == _GEN_8509 ? $signed(regsA_79_re) : $signed(_GEN_1142); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1144 = 8'h96 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1143); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1145 = 8'h97 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1144); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1146 = 8'h98 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1145); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1147 = 8'h99 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1146); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1148 = 8'h9a == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1147); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1149 = 8'h9b == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1148); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1150 = 8'h9c == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1149); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1151 = 8'h9d == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1150); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1152 = 8'h9e == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1151); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1153 = 8'h9f == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1152); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1154 = 8'ha0 == _GEN_8509 ? $signed(regsA_80_re) : $signed(_GEN_1153); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1155 = 8'ha1 == _GEN_8509 ? $signed(regsA_81_re) : $signed(_GEN_1154); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1156 = 8'ha2 == _GEN_8509 ? $signed(regsA_82_re) : $signed(_GEN_1155); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1157 = 8'ha3 == _GEN_8509 ? $signed(regsA_83_re) : $signed(_GEN_1156); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1158 = 8'ha4 == _GEN_8509 ? $signed(regsA_84_re) : $signed(_GEN_1157); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1159 = 8'ha5 == _GEN_8509 ? $signed(regsA_85_re) : $signed(_GEN_1158); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1160 = 8'ha6 == _GEN_8509 ? $signed(regsA_86_re) : $signed(_GEN_1159); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1161 = 8'ha7 == _GEN_8509 ? $signed(regsA_87_re) : $signed(_GEN_1160); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1162 = 8'ha8 == _GEN_8509 ? $signed(regsA_88_re) : $signed(_GEN_1161); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1163 = 8'ha9 == _GEN_8509 ? $signed(regsA_89_re) : $signed(_GEN_1162); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1164 = 8'haa == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1163); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1165 = 8'hab == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1164); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1166 = 8'hac == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1165); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1167 = 8'had == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1166); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1168 = 8'hae == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1167); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1169 = 8'haf == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1168); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1170 = 8'hb0 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1169); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1171 = 8'hb1 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1170); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1172 = 8'hb2 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1171); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1173 = 8'hb3 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_1172); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1174 = 8'hb4 == _GEN_8509 ? $signed(regsA_90_re) : $signed(_GEN_1173); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1175 = 8'hb5 == _GEN_8509 ? $signed(regsA_91_re) : $signed(_GEN_1174); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1176 = 8'hb6 == _GEN_8509 ? $signed(regsA_92_re) : $signed(_GEN_1175); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1177 = 8'hb7 == _GEN_8509 ? $signed(regsA_93_re) : $signed(_GEN_1176); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1178 = 8'hb8 == _GEN_8509 ? $signed(regsA_94_re) : $signed(_GEN_1177); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1179 = 8'hb9 == _GEN_8509 ? $signed(regsA_95_re) : $signed(_GEN_1178); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1180 = 8'hba == _GEN_8509 ? $signed(regsA_96_re) : $signed(_GEN_1179); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1181 = 8'hbb == _GEN_8509 ? $signed(regsA_97_re) : $signed(_GEN_1180); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1182 = 8'hbc == _GEN_8509 ? $signed(regsA_98_re) : $signed(_GEN_1181); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1183 = 8'hbd == _GEN_8509 ? $signed(regsA_99_re) : $signed(_GEN_1182); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [5:0] _T_4 = 1'h1 * 5'h13; // @[Matrix_Mul_V1.scala 148:44]
  wire [5:0] _T_6 = _T_4 + input_point; // @[Matrix_Mul_V1.scala 148:60]
  wire [31:0] _GEN_1185 = 6'h1 == _T_6 ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1186 = 6'h2 == _T_6 ? $signed(regsA_2_im) : $signed(_GEN_1185); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1187 = 6'h3 == _T_6 ? $signed(regsA_3_im) : $signed(_GEN_1186); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1188 = 6'h4 == _T_6 ? $signed(regsA_4_im) : $signed(_GEN_1187); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1189 = 6'h5 == _T_6 ? $signed(regsA_5_im) : $signed(_GEN_1188); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1190 = 6'h6 == _T_6 ? $signed(regsA_6_im) : $signed(_GEN_1189); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1191 = 6'h7 == _T_6 ? $signed(regsA_7_im) : $signed(_GEN_1190); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1192 = 6'h8 == _T_6 ? $signed(regsA_8_im) : $signed(_GEN_1191); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1193 = 6'h9 == _T_6 ? $signed(regsA_9_im) : $signed(_GEN_1192); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1194 = 6'ha == _T_6 ? $signed(32'sh0) : $signed(_GEN_1193); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1195 = 6'hb == _T_6 ? $signed(32'sh0) : $signed(_GEN_1194); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1196 = 6'hc == _T_6 ? $signed(32'sh0) : $signed(_GEN_1195); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1197 = 6'hd == _T_6 ? $signed(32'sh0) : $signed(_GEN_1196); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1198 = 6'he == _T_6 ? $signed(32'sh0) : $signed(_GEN_1197); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1199 = 6'hf == _T_6 ? $signed(32'sh0) : $signed(_GEN_1198); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1200 = 6'h10 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1199); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1201 = 6'h11 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1200); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1202 = 6'h12 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1201); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1203 = 6'h13 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1202); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1204 = 6'h14 == _T_6 ? $signed(regsA_10_im) : $signed(_GEN_1203); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1205 = 6'h15 == _T_6 ? $signed(regsA_11_im) : $signed(_GEN_1204); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1206 = 6'h16 == _T_6 ? $signed(regsA_12_im) : $signed(_GEN_1205); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1207 = 6'h17 == _T_6 ? $signed(regsA_13_im) : $signed(_GEN_1206); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1208 = 6'h18 == _T_6 ? $signed(regsA_14_im) : $signed(_GEN_1207); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1209 = 6'h19 == _T_6 ? $signed(regsA_15_im) : $signed(_GEN_1208); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1210 = 6'h1a == _T_6 ? $signed(regsA_16_im) : $signed(_GEN_1209); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1211 = 6'h1b == _T_6 ? $signed(regsA_17_im) : $signed(_GEN_1210); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1212 = 6'h1c == _T_6 ? $signed(regsA_18_im) : $signed(_GEN_1211); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1213 = 6'h1d == _T_6 ? $signed(regsA_19_im) : $signed(_GEN_1212); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1214 = 6'h1e == _T_6 ? $signed(32'sh0) : $signed(_GEN_1213); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1215 = 6'h1f == _T_6 ? $signed(32'sh0) : $signed(_GEN_1214); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1216 = 6'h20 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1215); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1217 = 6'h21 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1216); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1218 = 6'h22 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1217); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1219 = 6'h23 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1218); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1220 = 6'h24 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1219); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1221 = 6'h25 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1220); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1222 = 6'h26 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1221); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1223 = 6'h27 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1222); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1224 = 6'h28 == _T_6 ? $signed(regsA_20_im) : $signed(_GEN_1223); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1225 = 6'h29 == _T_6 ? $signed(regsA_21_im) : $signed(_GEN_1224); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1226 = 6'h2a == _T_6 ? $signed(regsA_22_im) : $signed(_GEN_1225); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1227 = 6'h2b == _T_6 ? $signed(regsA_23_im) : $signed(_GEN_1226); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1228 = 6'h2c == _T_6 ? $signed(regsA_24_im) : $signed(_GEN_1227); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1229 = 6'h2d == _T_6 ? $signed(regsA_25_im) : $signed(_GEN_1228); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1230 = 6'h2e == _T_6 ? $signed(regsA_26_im) : $signed(_GEN_1229); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1231 = 6'h2f == _T_6 ? $signed(regsA_27_im) : $signed(_GEN_1230); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1232 = 6'h30 == _T_6 ? $signed(regsA_28_im) : $signed(_GEN_1231); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1233 = 6'h31 == _T_6 ? $signed(regsA_29_im) : $signed(_GEN_1232); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1234 = 6'h32 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1233); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1235 = 6'h33 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1234); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1236 = 6'h34 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1235); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1237 = 6'h35 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1236); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1238 = 6'h36 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1237); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1239 = 6'h37 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1238); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1240 = 6'h38 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1239); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1241 = 6'h39 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1240); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1242 = 6'h3a == _T_6 ? $signed(32'sh0) : $signed(_GEN_1241); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1243 = 6'h3b == _T_6 ? $signed(32'sh0) : $signed(_GEN_1242); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1244 = 6'h3c == _T_6 ? $signed(regsA_30_im) : $signed(_GEN_1243); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1245 = 6'h3d == _T_6 ? $signed(regsA_31_im) : $signed(_GEN_1244); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1246 = 6'h3e == _T_6 ? $signed(regsA_32_im) : $signed(_GEN_1245); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1247 = 6'h3f == _T_6 ? $signed(regsA_33_im) : $signed(_GEN_1246); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [6:0] _GEN_8697 = {{1'd0}, _T_6}; // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1248 = 7'h40 == _GEN_8697 ? $signed(regsA_34_im) : $signed(_GEN_1247); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1249 = 7'h41 == _GEN_8697 ? $signed(regsA_35_im) : $signed(_GEN_1248); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1250 = 7'h42 == _GEN_8697 ? $signed(regsA_36_im) : $signed(_GEN_1249); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1251 = 7'h43 == _GEN_8697 ? $signed(regsA_37_im) : $signed(_GEN_1250); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1252 = 7'h44 == _GEN_8697 ? $signed(regsA_38_im) : $signed(_GEN_1251); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1253 = 7'h45 == _GEN_8697 ? $signed(regsA_39_im) : $signed(_GEN_1252); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1254 = 7'h46 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1253); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1255 = 7'h47 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1254); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1256 = 7'h48 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1255); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1257 = 7'h49 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1256); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1258 = 7'h4a == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1257); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1259 = 7'h4b == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1258); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1260 = 7'h4c == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1259); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1261 = 7'h4d == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1260); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1262 = 7'h4e == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1261); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1263 = 7'h4f == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1262); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1264 = 7'h50 == _GEN_8697 ? $signed(regsA_40_im) : $signed(_GEN_1263); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1265 = 7'h51 == _GEN_8697 ? $signed(regsA_41_im) : $signed(_GEN_1264); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1266 = 7'h52 == _GEN_8697 ? $signed(regsA_42_im) : $signed(_GEN_1265); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1267 = 7'h53 == _GEN_8697 ? $signed(regsA_43_im) : $signed(_GEN_1266); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1268 = 7'h54 == _GEN_8697 ? $signed(regsA_44_im) : $signed(_GEN_1267); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1269 = 7'h55 == _GEN_8697 ? $signed(regsA_45_im) : $signed(_GEN_1268); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1270 = 7'h56 == _GEN_8697 ? $signed(regsA_46_im) : $signed(_GEN_1269); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1271 = 7'h57 == _GEN_8697 ? $signed(regsA_47_im) : $signed(_GEN_1270); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1272 = 7'h58 == _GEN_8697 ? $signed(regsA_48_im) : $signed(_GEN_1271); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1273 = 7'h59 == _GEN_8697 ? $signed(regsA_49_im) : $signed(_GEN_1272); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1274 = 7'h5a == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1273); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1275 = 7'h5b == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1274); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1276 = 7'h5c == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1275); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1277 = 7'h5d == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1276); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1278 = 7'h5e == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1277); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1279 = 7'h5f == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1278); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1280 = 7'h60 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1279); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1281 = 7'h61 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1280); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1282 = 7'h62 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1281); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1283 = 7'h63 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1282); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1284 = 7'h64 == _GEN_8697 ? $signed(regsA_50_im) : $signed(_GEN_1283); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1285 = 7'h65 == _GEN_8697 ? $signed(regsA_51_im) : $signed(_GEN_1284); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1286 = 7'h66 == _GEN_8697 ? $signed(regsA_52_im) : $signed(_GEN_1285); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1287 = 7'h67 == _GEN_8697 ? $signed(regsA_53_im) : $signed(_GEN_1286); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1288 = 7'h68 == _GEN_8697 ? $signed(regsA_54_im) : $signed(_GEN_1287); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1289 = 7'h69 == _GEN_8697 ? $signed(regsA_55_im) : $signed(_GEN_1288); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1290 = 7'h6a == _GEN_8697 ? $signed(regsA_56_im) : $signed(_GEN_1289); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1291 = 7'h6b == _GEN_8697 ? $signed(regsA_57_im) : $signed(_GEN_1290); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1292 = 7'h6c == _GEN_8697 ? $signed(regsA_58_im) : $signed(_GEN_1291); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1293 = 7'h6d == _GEN_8697 ? $signed(regsA_59_im) : $signed(_GEN_1292); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1294 = 7'h6e == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1293); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1295 = 7'h6f == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1294); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1296 = 7'h70 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1295); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1297 = 7'h71 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1296); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1298 = 7'h72 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1297); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1299 = 7'h73 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1298); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1300 = 7'h74 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1299); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1301 = 7'h75 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1300); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1302 = 7'h76 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1301); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1303 = 7'h77 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1302); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1304 = 7'h78 == _GEN_8697 ? $signed(regsA_60_im) : $signed(_GEN_1303); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1305 = 7'h79 == _GEN_8697 ? $signed(regsA_61_im) : $signed(_GEN_1304); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1306 = 7'h7a == _GEN_8697 ? $signed(regsA_62_im) : $signed(_GEN_1305); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1307 = 7'h7b == _GEN_8697 ? $signed(regsA_63_im) : $signed(_GEN_1306); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1308 = 7'h7c == _GEN_8697 ? $signed(regsA_64_im) : $signed(_GEN_1307); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1309 = 7'h7d == _GEN_8697 ? $signed(regsA_65_im) : $signed(_GEN_1308); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1310 = 7'h7e == _GEN_8697 ? $signed(regsA_66_im) : $signed(_GEN_1309); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1311 = 7'h7f == _GEN_8697 ? $signed(regsA_67_im) : $signed(_GEN_1310); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [7:0] _GEN_8761 = {{2'd0}, _T_6}; // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1312 = 8'h80 == _GEN_8761 ? $signed(regsA_68_im) : $signed(_GEN_1311); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1313 = 8'h81 == _GEN_8761 ? $signed(regsA_69_im) : $signed(_GEN_1312); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1314 = 8'h82 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1313); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1315 = 8'h83 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1314); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1316 = 8'h84 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1315); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1317 = 8'h85 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1316); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1318 = 8'h86 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1317); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1319 = 8'h87 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1318); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1320 = 8'h88 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1319); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1321 = 8'h89 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1320); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1322 = 8'h8a == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1321); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1323 = 8'h8b == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1322); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1324 = 8'h8c == _GEN_8761 ? $signed(regsA_70_im) : $signed(_GEN_1323); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1325 = 8'h8d == _GEN_8761 ? $signed(regsA_71_im) : $signed(_GEN_1324); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1326 = 8'h8e == _GEN_8761 ? $signed(regsA_72_im) : $signed(_GEN_1325); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1327 = 8'h8f == _GEN_8761 ? $signed(regsA_73_im) : $signed(_GEN_1326); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1328 = 8'h90 == _GEN_8761 ? $signed(regsA_74_im) : $signed(_GEN_1327); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1329 = 8'h91 == _GEN_8761 ? $signed(regsA_75_im) : $signed(_GEN_1328); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1330 = 8'h92 == _GEN_8761 ? $signed(regsA_76_im) : $signed(_GEN_1329); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1331 = 8'h93 == _GEN_8761 ? $signed(regsA_77_im) : $signed(_GEN_1330); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1332 = 8'h94 == _GEN_8761 ? $signed(regsA_78_im) : $signed(_GEN_1331); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1333 = 8'h95 == _GEN_8761 ? $signed(regsA_79_im) : $signed(_GEN_1332); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1334 = 8'h96 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1333); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1335 = 8'h97 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1334); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1336 = 8'h98 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1335); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1337 = 8'h99 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1336); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1338 = 8'h9a == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1337); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1339 = 8'h9b == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1338); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1340 = 8'h9c == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1339); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1341 = 8'h9d == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1340); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1342 = 8'h9e == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1341); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1343 = 8'h9f == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1342); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1344 = 8'ha0 == _GEN_8761 ? $signed(regsA_80_im) : $signed(_GEN_1343); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1345 = 8'ha1 == _GEN_8761 ? $signed(regsA_81_im) : $signed(_GEN_1344); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1346 = 8'ha2 == _GEN_8761 ? $signed(regsA_82_im) : $signed(_GEN_1345); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1347 = 8'ha3 == _GEN_8761 ? $signed(regsA_83_im) : $signed(_GEN_1346); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1348 = 8'ha4 == _GEN_8761 ? $signed(regsA_84_im) : $signed(_GEN_1347); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1349 = 8'ha5 == _GEN_8761 ? $signed(regsA_85_im) : $signed(_GEN_1348); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1350 = 8'ha6 == _GEN_8761 ? $signed(regsA_86_im) : $signed(_GEN_1349); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1351 = 8'ha7 == _GEN_8761 ? $signed(regsA_87_im) : $signed(_GEN_1350); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1352 = 8'ha8 == _GEN_8761 ? $signed(regsA_88_im) : $signed(_GEN_1351); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1353 = 8'ha9 == _GEN_8761 ? $signed(regsA_89_im) : $signed(_GEN_1352); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1354 = 8'haa == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1353); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1355 = 8'hab == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1354); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1356 = 8'hac == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1355); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1357 = 8'had == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1356); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1358 = 8'hae == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1357); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1359 = 8'haf == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1358); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1360 = 8'hb0 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1359); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1361 = 8'hb1 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1360); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1362 = 8'hb2 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1361); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1363 = 8'hb3 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1362); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1364 = 8'hb4 == _GEN_8761 ? $signed(regsA_90_im) : $signed(_GEN_1363); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1365 = 8'hb5 == _GEN_8761 ? $signed(regsA_91_im) : $signed(_GEN_1364); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1366 = 8'hb6 == _GEN_8761 ? $signed(regsA_92_im) : $signed(_GEN_1365); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1367 = 8'hb7 == _GEN_8761 ? $signed(regsA_93_im) : $signed(_GEN_1366); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1368 = 8'hb8 == _GEN_8761 ? $signed(regsA_94_im) : $signed(_GEN_1367); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1369 = 8'hb9 == _GEN_8761 ? $signed(regsA_95_im) : $signed(_GEN_1368); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1370 = 8'hba == _GEN_8761 ? $signed(regsA_96_im) : $signed(_GEN_1369); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1371 = 8'hbb == _GEN_8761 ? $signed(regsA_97_im) : $signed(_GEN_1370); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1372 = 8'hbc == _GEN_8761 ? $signed(regsA_98_im) : $signed(_GEN_1371); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1373 = 8'hbd == _GEN_8761 ? $signed(regsA_99_im) : $signed(_GEN_1372); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1375 = 6'h1 == _T_6 ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1376 = 6'h2 == _T_6 ? $signed(regsA_2_re) : $signed(_GEN_1375); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1377 = 6'h3 == _T_6 ? $signed(regsA_3_re) : $signed(_GEN_1376); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1378 = 6'h4 == _T_6 ? $signed(regsA_4_re) : $signed(_GEN_1377); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1379 = 6'h5 == _T_6 ? $signed(regsA_5_re) : $signed(_GEN_1378); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1380 = 6'h6 == _T_6 ? $signed(regsA_6_re) : $signed(_GEN_1379); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1381 = 6'h7 == _T_6 ? $signed(regsA_7_re) : $signed(_GEN_1380); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1382 = 6'h8 == _T_6 ? $signed(regsA_8_re) : $signed(_GEN_1381); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1383 = 6'h9 == _T_6 ? $signed(regsA_9_re) : $signed(_GEN_1382); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1384 = 6'ha == _T_6 ? $signed(32'sh0) : $signed(_GEN_1383); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1385 = 6'hb == _T_6 ? $signed(32'sh0) : $signed(_GEN_1384); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1386 = 6'hc == _T_6 ? $signed(32'sh0) : $signed(_GEN_1385); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1387 = 6'hd == _T_6 ? $signed(32'sh0) : $signed(_GEN_1386); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1388 = 6'he == _T_6 ? $signed(32'sh0) : $signed(_GEN_1387); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1389 = 6'hf == _T_6 ? $signed(32'sh0) : $signed(_GEN_1388); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1390 = 6'h10 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1389); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1391 = 6'h11 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1390); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1392 = 6'h12 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1391); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1393 = 6'h13 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1392); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1394 = 6'h14 == _T_6 ? $signed(regsA_10_re) : $signed(_GEN_1393); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1395 = 6'h15 == _T_6 ? $signed(regsA_11_re) : $signed(_GEN_1394); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1396 = 6'h16 == _T_6 ? $signed(regsA_12_re) : $signed(_GEN_1395); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1397 = 6'h17 == _T_6 ? $signed(regsA_13_re) : $signed(_GEN_1396); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1398 = 6'h18 == _T_6 ? $signed(regsA_14_re) : $signed(_GEN_1397); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1399 = 6'h19 == _T_6 ? $signed(regsA_15_re) : $signed(_GEN_1398); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1400 = 6'h1a == _T_6 ? $signed(regsA_16_re) : $signed(_GEN_1399); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1401 = 6'h1b == _T_6 ? $signed(regsA_17_re) : $signed(_GEN_1400); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1402 = 6'h1c == _T_6 ? $signed(regsA_18_re) : $signed(_GEN_1401); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1403 = 6'h1d == _T_6 ? $signed(regsA_19_re) : $signed(_GEN_1402); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1404 = 6'h1e == _T_6 ? $signed(32'sh0) : $signed(_GEN_1403); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1405 = 6'h1f == _T_6 ? $signed(32'sh0) : $signed(_GEN_1404); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1406 = 6'h20 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1405); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1407 = 6'h21 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1406); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1408 = 6'h22 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1407); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1409 = 6'h23 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1408); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1410 = 6'h24 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1409); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1411 = 6'h25 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1410); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1412 = 6'h26 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1411); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1413 = 6'h27 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1412); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1414 = 6'h28 == _T_6 ? $signed(regsA_20_re) : $signed(_GEN_1413); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1415 = 6'h29 == _T_6 ? $signed(regsA_21_re) : $signed(_GEN_1414); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1416 = 6'h2a == _T_6 ? $signed(regsA_22_re) : $signed(_GEN_1415); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1417 = 6'h2b == _T_6 ? $signed(regsA_23_re) : $signed(_GEN_1416); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1418 = 6'h2c == _T_6 ? $signed(regsA_24_re) : $signed(_GEN_1417); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1419 = 6'h2d == _T_6 ? $signed(regsA_25_re) : $signed(_GEN_1418); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1420 = 6'h2e == _T_6 ? $signed(regsA_26_re) : $signed(_GEN_1419); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1421 = 6'h2f == _T_6 ? $signed(regsA_27_re) : $signed(_GEN_1420); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1422 = 6'h30 == _T_6 ? $signed(regsA_28_re) : $signed(_GEN_1421); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1423 = 6'h31 == _T_6 ? $signed(regsA_29_re) : $signed(_GEN_1422); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1424 = 6'h32 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1423); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1425 = 6'h33 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1424); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1426 = 6'h34 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1425); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1427 = 6'h35 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1426); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1428 = 6'h36 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1427); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1429 = 6'h37 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1428); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1430 = 6'h38 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1429); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1431 = 6'h39 == _T_6 ? $signed(32'sh0) : $signed(_GEN_1430); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1432 = 6'h3a == _T_6 ? $signed(32'sh0) : $signed(_GEN_1431); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1433 = 6'h3b == _T_6 ? $signed(32'sh0) : $signed(_GEN_1432); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1434 = 6'h3c == _T_6 ? $signed(regsA_30_re) : $signed(_GEN_1433); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1435 = 6'h3d == _T_6 ? $signed(regsA_31_re) : $signed(_GEN_1434); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1436 = 6'h3e == _T_6 ? $signed(regsA_32_re) : $signed(_GEN_1435); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1437 = 6'h3f == _T_6 ? $signed(regsA_33_re) : $signed(_GEN_1436); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1438 = 7'h40 == _GEN_8697 ? $signed(regsA_34_re) : $signed(_GEN_1437); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1439 = 7'h41 == _GEN_8697 ? $signed(regsA_35_re) : $signed(_GEN_1438); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1440 = 7'h42 == _GEN_8697 ? $signed(regsA_36_re) : $signed(_GEN_1439); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1441 = 7'h43 == _GEN_8697 ? $signed(regsA_37_re) : $signed(_GEN_1440); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1442 = 7'h44 == _GEN_8697 ? $signed(regsA_38_re) : $signed(_GEN_1441); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1443 = 7'h45 == _GEN_8697 ? $signed(regsA_39_re) : $signed(_GEN_1442); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1444 = 7'h46 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1443); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1445 = 7'h47 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1444); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1446 = 7'h48 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1445); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1447 = 7'h49 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1446); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1448 = 7'h4a == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1447); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1449 = 7'h4b == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1448); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1450 = 7'h4c == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1449); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1451 = 7'h4d == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1450); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1452 = 7'h4e == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1451); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1453 = 7'h4f == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1452); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1454 = 7'h50 == _GEN_8697 ? $signed(regsA_40_re) : $signed(_GEN_1453); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1455 = 7'h51 == _GEN_8697 ? $signed(regsA_41_re) : $signed(_GEN_1454); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1456 = 7'h52 == _GEN_8697 ? $signed(regsA_42_re) : $signed(_GEN_1455); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1457 = 7'h53 == _GEN_8697 ? $signed(regsA_43_re) : $signed(_GEN_1456); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1458 = 7'h54 == _GEN_8697 ? $signed(regsA_44_re) : $signed(_GEN_1457); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1459 = 7'h55 == _GEN_8697 ? $signed(regsA_45_re) : $signed(_GEN_1458); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1460 = 7'h56 == _GEN_8697 ? $signed(regsA_46_re) : $signed(_GEN_1459); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1461 = 7'h57 == _GEN_8697 ? $signed(regsA_47_re) : $signed(_GEN_1460); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1462 = 7'h58 == _GEN_8697 ? $signed(regsA_48_re) : $signed(_GEN_1461); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1463 = 7'h59 == _GEN_8697 ? $signed(regsA_49_re) : $signed(_GEN_1462); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1464 = 7'h5a == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1463); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1465 = 7'h5b == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1464); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1466 = 7'h5c == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1465); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1467 = 7'h5d == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1466); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1468 = 7'h5e == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1467); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1469 = 7'h5f == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1468); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1470 = 7'h60 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1469); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1471 = 7'h61 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1470); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1472 = 7'h62 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1471); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1473 = 7'h63 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1472); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1474 = 7'h64 == _GEN_8697 ? $signed(regsA_50_re) : $signed(_GEN_1473); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1475 = 7'h65 == _GEN_8697 ? $signed(regsA_51_re) : $signed(_GEN_1474); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1476 = 7'h66 == _GEN_8697 ? $signed(regsA_52_re) : $signed(_GEN_1475); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1477 = 7'h67 == _GEN_8697 ? $signed(regsA_53_re) : $signed(_GEN_1476); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1478 = 7'h68 == _GEN_8697 ? $signed(regsA_54_re) : $signed(_GEN_1477); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1479 = 7'h69 == _GEN_8697 ? $signed(regsA_55_re) : $signed(_GEN_1478); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1480 = 7'h6a == _GEN_8697 ? $signed(regsA_56_re) : $signed(_GEN_1479); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1481 = 7'h6b == _GEN_8697 ? $signed(regsA_57_re) : $signed(_GEN_1480); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1482 = 7'h6c == _GEN_8697 ? $signed(regsA_58_re) : $signed(_GEN_1481); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1483 = 7'h6d == _GEN_8697 ? $signed(regsA_59_re) : $signed(_GEN_1482); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1484 = 7'h6e == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1483); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1485 = 7'h6f == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1484); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1486 = 7'h70 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1485); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1487 = 7'h71 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1486); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1488 = 7'h72 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1487); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1489 = 7'h73 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1488); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1490 = 7'h74 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1489); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1491 = 7'h75 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1490); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1492 = 7'h76 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1491); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1493 = 7'h77 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_1492); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1494 = 7'h78 == _GEN_8697 ? $signed(regsA_60_re) : $signed(_GEN_1493); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1495 = 7'h79 == _GEN_8697 ? $signed(regsA_61_re) : $signed(_GEN_1494); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1496 = 7'h7a == _GEN_8697 ? $signed(regsA_62_re) : $signed(_GEN_1495); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1497 = 7'h7b == _GEN_8697 ? $signed(regsA_63_re) : $signed(_GEN_1496); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1498 = 7'h7c == _GEN_8697 ? $signed(regsA_64_re) : $signed(_GEN_1497); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1499 = 7'h7d == _GEN_8697 ? $signed(regsA_65_re) : $signed(_GEN_1498); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1500 = 7'h7e == _GEN_8697 ? $signed(regsA_66_re) : $signed(_GEN_1499); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1501 = 7'h7f == _GEN_8697 ? $signed(regsA_67_re) : $signed(_GEN_1500); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1502 = 8'h80 == _GEN_8761 ? $signed(regsA_68_re) : $signed(_GEN_1501); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1503 = 8'h81 == _GEN_8761 ? $signed(regsA_69_re) : $signed(_GEN_1502); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1504 = 8'h82 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1503); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1505 = 8'h83 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1504); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1506 = 8'h84 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1505); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1507 = 8'h85 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1506); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1508 = 8'h86 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1507); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1509 = 8'h87 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1508); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1510 = 8'h88 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1509); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1511 = 8'h89 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1510); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1512 = 8'h8a == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1511); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1513 = 8'h8b == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1512); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1514 = 8'h8c == _GEN_8761 ? $signed(regsA_70_re) : $signed(_GEN_1513); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1515 = 8'h8d == _GEN_8761 ? $signed(regsA_71_re) : $signed(_GEN_1514); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1516 = 8'h8e == _GEN_8761 ? $signed(regsA_72_re) : $signed(_GEN_1515); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1517 = 8'h8f == _GEN_8761 ? $signed(regsA_73_re) : $signed(_GEN_1516); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1518 = 8'h90 == _GEN_8761 ? $signed(regsA_74_re) : $signed(_GEN_1517); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1519 = 8'h91 == _GEN_8761 ? $signed(regsA_75_re) : $signed(_GEN_1518); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1520 = 8'h92 == _GEN_8761 ? $signed(regsA_76_re) : $signed(_GEN_1519); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1521 = 8'h93 == _GEN_8761 ? $signed(regsA_77_re) : $signed(_GEN_1520); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1522 = 8'h94 == _GEN_8761 ? $signed(regsA_78_re) : $signed(_GEN_1521); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1523 = 8'h95 == _GEN_8761 ? $signed(regsA_79_re) : $signed(_GEN_1522); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1524 = 8'h96 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1523); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1525 = 8'h97 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1524); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1526 = 8'h98 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1525); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1527 = 8'h99 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1526); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1528 = 8'h9a == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1527); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1529 = 8'h9b == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1528); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1530 = 8'h9c == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1529); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1531 = 8'h9d == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1530); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1532 = 8'h9e == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1531); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1533 = 8'h9f == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1532); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1534 = 8'ha0 == _GEN_8761 ? $signed(regsA_80_re) : $signed(_GEN_1533); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1535 = 8'ha1 == _GEN_8761 ? $signed(regsA_81_re) : $signed(_GEN_1534); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1536 = 8'ha2 == _GEN_8761 ? $signed(regsA_82_re) : $signed(_GEN_1535); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1537 = 8'ha3 == _GEN_8761 ? $signed(regsA_83_re) : $signed(_GEN_1536); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1538 = 8'ha4 == _GEN_8761 ? $signed(regsA_84_re) : $signed(_GEN_1537); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1539 = 8'ha5 == _GEN_8761 ? $signed(regsA_85_re) : $signed(_GEN_1538); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1540 = 8'ha6 == _GEN_8761 ? $signed(regsA_86_re) : $signed(_GEN_1539); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1541 = 8'ha7 == _GEN_8761 ? $signed(regsA_87_re) : $signed(_GEN_1540); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1542 = 8'ha8 == _GEN_8761 ? $signed(regsA_88_re) : $signed(_GEN_1541); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1543 = 8'ha9 == _GEN_8761 ? $signed(regsA_89_re) : $signed(_GEN_1542); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1544 = 8'haa == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1543); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1545 = 8'hab == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1544); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1546 = 8'hac == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1545); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1547 = 8'had == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1546); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1548 = 8'hae == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1547); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1549 = 8'haf == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1548); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1550 = 8'hb0 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1549); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1551 = 8'hb1 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1550); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1552 = 8'hb2 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1551); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1553 = 8'hb3 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_1552); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1554 = 8'hb4 == _GEN_8761 ? $signed(regsA_90_re) : $signed(_GEN_1553); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1555 = 8'hb5 == _GEN_8761 ? $signed(regsA_91_re) : $signed(_GEN_1554); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1556 = 8'hb6 == _GEN_8761 ? $signed(regsA_92_re) : $signed(_GEN_1555); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1557 = 8'hb7 == _GEN_8761 ? $signed(regsA_93_re) : $signed(_GEN_1556); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1558 = 8'hb8 == _GEN_8761 ? $signed(regsA_94_re) : $signed(_GEN_1557); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1559 = 8'hb9 == _GEN_8761 ? $signed(regsA_95_re) : $signed(_GEN_1558); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1560 = 8'hba == _GEN_8761 ? $signed(regsA_96_re) : $signed(_GEN_1559); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1561 = 8'hbb == _GEN_8761 ? $signed(regsA_97_re) : $signed(_GEN_1560); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1562 = 8'hbc == _GEN_8761 ? $signed(regsA_98_re) : $signed(_GEN_1561); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1563 = 8'hbd == _GEN_8761 ? $signed(regsA_99_re) : $signed(_GEN_1562); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [6:0] _T_7 = 2'h2 * 5'h13; // @[Matrix_Mul_V1.scala 148:44]
  wire [6:0] _GEN_8949 = {{1'd0}, input_point}; // @[Matrix_Mul_V1.scala 148:60]
  wire [6:0] _T_9 = _T_7 + _GEN_8949; // @[Matrix_Mul_V1.scala 148:60]
  wire [31:0] _GEN_1565 = 7'h1 == _T_9 ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1566 = 7'h2 == _T_9 ? $signed(regsA_2_im) : $signed(_GEN_1565); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1567 = 7'h3 == _T_9 ? $signed(regsA_3_im) : $signed(_GEN_1566); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1568 = 7'h4 == _T_9 ? $signed(regsA_4_im) : $signed(_GEN_1567); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1569 = 7'h5 == _T_9 ? $signed(regsA_5_im) : $signed(_GEN_1568); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1570 = 7'h6 == _T_9 ? $signed(regsA_6_im) : $signed(_GEN_1569); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1571 = 7'h7 == _T_9 ? $signed(regsA_7_im) : $signed(_GEN_1570); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1572 = 7'h8 == _T_9 ? $signed(regsA_8_im) : $signed(_GEN_1571); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1573 = 7'h9 == _T_9 ? $signed(regsA_9_im) : $signed(_GEN_1572); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1574 = 7'ha == _T_9 ? $signed(32'sh0) : $signed(_GEN_1573); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1575 = 7'hb == _T_9 ? $signed(32'sh0) : $signed(_GEN_1574); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1576 = 7'hc == _T_9 ? $signed(32'sh0) : $signed(_GEN_1575); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1577 = 7'hd == _T_9 ? $signed(32'sh0) : $signed(_GEN_1576); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1578 = 7'he == _T_9 ? $signed(32'sh0) : $signed(_GEN_1577); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1579 = 7'hf == _T_9 ? $signed(32'sh0) : $signed(_GEN_1578); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1580 = 7'h10 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1579); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1581 = 7'h11 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1580); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1582 = 7'h12 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1581); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1583 = 7'h13 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1582); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1584 = 7'h14 == _T_9 ? $signed(regsA_10_im) : $signed(_GEN_1583); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1585 = 7'h15 == _T_9 ? $signed(regsA_11_im) : $signed(_GEN_1584); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1586 = 7'h16 == _T_9 ? $signed(regsA_12_im) : $signed(_GEN_1585); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1587 = 7'h17 == _T_9 ? $signed(regsA_13_im) : $signed(_GEN_1586); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1588 = 7'h18 == _T_9 ? $signed(regsA_14_im) : $signed(_GEN_1587); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1589 = 7'h19 == _T_9 ? $signed(regsA_15_im) : $signed(_GEN_1588); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1590 = 7'h1a == _T_9 ? $signed(regsA_16_im) : $signed(_GEN_1589); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1591 = 7'h1b == _T_9 ? $signed(regsA_17_im) : $signed(_GEN_1590); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1592 = 7'h1c == _T_9 ? $signed(regsA_18_im) : $signed(_GEN_1591); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1593 = 7'h1d == _T_9 ? $signed(regsA_19_im) : $signed(_GEN_1592); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1594 = 7'h1e == _T_9 ? $signed(32'sh0) : $signed(_GEN_1593); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1595 = 7'h1f == _T_9 ? $signed(32'sh0) : $signed(_GEN_1594); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1596 = 7'h20 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1595); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1597 = 7'h21 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1596); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1598 = 7'h22 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1597); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1599 = 7'h23 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1598); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1600 = 7'h24 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1599); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1601 = 7'h25 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1600); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1602 = 7'h26 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1601); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1603 = 7'h27 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1602); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1604 = 7'h28 == _T_9 ? $signed(regsA_20_im) : $signed(_GEN_1603); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1605 = 7'h29 == _T_9 ? $signed(regsA_21_im) : $signed(_GEN_1604); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1606 = 7'h2a == _T_9 ? $signed(regsA_22_im) : $signed(_GEN_1605); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1607 = 7'h2b == _T_9 ? $signed(regsA_23_im) : $signed(_GEN_1606); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1608 = 7'h2c == _T_9 ? $signed(regsA_24_im) : $signed(_GEN_1607); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1609 = 7'h2d == _T_9 ? $signed(regsA_25_im) : $signed(_GEN_1608); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1610 = 7'h2e == _T_9 ? $signed(regsA_26_im) : $signed(_GEN_1609); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1611 = 7'h2f == _T_9 ? $signed(regsA_27_im) : $signed(_GEN_1610); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1612 = 7'h30 == _T_9 ? $signed(regsA_28_im) : $signed(_GEN_1611); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1613 = 7'h31 == _T_9 ? $signed(regsA_29_im) : $signed(_GEN_1612); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1614 = 7'h32 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1613); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1615 = 7'h33 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1614); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1616 = 7'h34 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1615); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1617 = 7'h35 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1616); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1618 = 7'h36 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1617); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1619 = 7'h37 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1618); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1620 = 7'h38 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1619); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1621 = 7'h39 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1620); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1622 = 7'h3a == _T_9 ? $signed(32'sh0) : $signed(_GEN_1621); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1623 = 7'h3b == _T_9 ? $signed(32'sh0) : $signed(_GEN_1622); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1624 = 7'h3c == _T_9 ? $signed(regsA_30_im) : $signed(_GEN_1623); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1625 = 7'h3d == _T_9 ? $signed(regsA_31_im) : $signed(_GEN_1624); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1626 = 7'h3e == _T_9 ? $signed(regsA_32_im) : $signed(_GEN_1625); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1627 = 7'h3f == _T_9 ? $signed(regsA_33_im) : $signed(_GEN_1626); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1628 = 7'h40 == _T_9 ? $signed(regsA_34_im) : $signed(_GEN_1627); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1629 = 7'h41 == _T_9 ? $signed(regsA_35_im) : $signed(_GEN_1628); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1630 = 7'h42 == _T_9 ? $signed(regsA_36_im) : $signed(_GEN_1629); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1631 = 7'h43 == _T_9 ? $signed(regsA_37_im) : $signed(_GEN_1630); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1632 = 7'h44 == _T_9 ? $signed(regsA_38_im) : $signed(_GEN_1631); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1633 = 7'h45 == _T_9 ? $signed(regsA_39_im) : $signed(_GEN_1632); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1634 = 7'h46 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1633); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1635 = 7'h47 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1634); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1636 = 7'h48 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1635); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1637 = 7'h49 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1636); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1638 = 7'h4a == _T_9 ? $signed(32'sh0) : $signed(_GEN_1637); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1639 = 7'h4b == _T_9 ? $signed(32'sh0) : $signed(_GEN_1638); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1640 = 7'h4c == _T_9 ? $signed(32'sh0) : $signed(_GEN_1639); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1641 = 7'h4d == _T_9 ? $signed(32'sh0) : $signed(_GEN_1640); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1642 = 7'h4e == _T_9 ? $signed(32'sh0) : $signed(_GEN_1641); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1643 = 7'h4f == _T_9 ? $signed(32'sh0) : $signed(_GEN_1642); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1644 = 7'h50 == _T_9 ? $signed(regsA_40_im) : $signed(_GEN_1643); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1645 = 7'h51 == _T_9 ? $signed(regsA_41_im) : $signed(_GEN_1644); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1646 = 7'h52 == _T_9 ? $signed(regsA_42_im) : $signed(_GEN_1645); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1647 = 7'h53 == _T_9 ? $signed(regsA_43_im) : $signed(_GEN_1646); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1648 = 7'h54 == _T_9 ? $signed(regsA_44_im) : $signed(_GEN_1647); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1649 = 7'h55 == _T_9 ? $signed(regsA_45_im) : $signed(_GEN_1648); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1650 = 7'h56 == _T_9 ? $signed(regsA_46_im) : $signed(_GEN_1649); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1651 = 7'h57 == _T_9 ? $signed(regsA_47_im) : $signed(_GEN_1650); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1652 = 7'h58 == _T_9 ? $signed(regsA_48_im) : $signed(_GEN_1651); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1653 = 7'h59 == _T_9 ? $signed(regsA_49_im) : $signed(_GEN_1652); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1654 = 7'h5a == _T_9 ? $signed(32'sh0) : $signed(_GEN_1653); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1655 = 7'h5b == _T_9 ? $signed(32'sh0) : $signed(_GEN_1654); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1656 = 7'h5c == _T_9 ? $signed(32'sh0) : $signed(_GEN_1655); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1657 = 7'h5d == _T_9 ? $signed(32'sh0) : $signed(_GEN_1656); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1658 = 7'h5e == _T_9 ? $signed(32'sh0) : $signed(_GEN_1657); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1659 = 7'h5f == _T_9 ? $signed(32'sh0) : $signed(_GEN_1658); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1660 = 7'h60 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1659); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1661 = 7'h61 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1660); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1662 = 7'h62 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1661); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1663 = 7'h63 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1662); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1664 = 7'h64 == _T_9 ? $signed(regsA_50_im) : $signed(_GEN_1663); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1665 = 7'h65 == _T_9 ? $signed(regsA_51_im) : $signed(_GEN_1664); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1666 = 7'h66 == _T_9 ? $signed(regsA_52_im) : $signed(_GEN_1665); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1667 = 7'h67 == _T_9 ? $signed(regsA_53_im) : $signed(_GEN_1666); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1668 = 7'h68 == _T_9 ? $signed(regsA_54_im) : $signed(_GEN_1667); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1669 = 7'h69 == _T_9 ? $signed(regsA_55_im) : $signed(_GEN_1668); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1670 = 7'h6a == _T_9 ? $signed(regsA_56_im) : $signed(_GEN_1669); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1671 = 7'h6b == _T_9 ? $signed(regsA_57_im) : $signed(_GEN_1670); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1672 = 7'h6c == _T_9 ? $signed(regsA_58_im) : $signed(_GEN_1671); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1673 = 7'h6d == _T_9 ? $signed(regsA_59_im) : $signed(_GEN_1672); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1674 = 7'h6e == _T_9 ? $signed(32'sh0) : $signed(_GEN_1673); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1675 = 7'h6f == _T_9 ? $signed(32'sh0) : $signed(_GEN_1674); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1676 = 7'h70 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1675); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1677 = 7'h71 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1676); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1678 = 7'h72 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1677); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1679 = 7'h73 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1678); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1680 = 7'h74 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1679); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1681 = 7'h75 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1680); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1682 = 7'h76 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1681); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1683 = 7'h77 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1682); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1684 = 7'h78 == _T_9 ? $signed(regsA_60_im) : $signed(_GEN_1683); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1685 = 7'h79 == _T_9 ? $signed(regsA_61_im) : $signed(_GEN_1684); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1686 = 7'h7a == _T_9 ? $signed(regsA_62_im) : $signed(_GEN_1685); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1687 = 7'h7b == _T_9 ? $signed(regsA_63_im) : $signed(_GEN_1686); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1688 = 7'h7c == _T_9 ? $signed(regsA_64_im) : $signed(_GEN_1687); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1689 = 7'h7d == _T_9 ? $signed(regsA_65_im) : $signed(_GEN_1688); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1690 = 7'h7e == _T_9 ? $signed(regsA_66_im) : $signed(_GEN_1689); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1691 = 7'h7f == _T_9 ? $signed(regsA_67_im) : $signed(_GEN_1690); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [7:0] _GEN_8950 = {{1'd0}, _T_9}; // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1692 = 8'h80 == _GEN_8950 ? $signed(regsA_68_im) : $signed(_GEN_1691); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1693 = 8'h81 == _GEN_8950 ? $signed(regsA_69_im) : $signed(_GEN_1692); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1694 = 8'h82 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1693); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1695 = 8'h83 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1694); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1696 = 8'h84 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1695); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1697 = 8'h85 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1696); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1698 = 8'h86 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1697); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1699 = 8'h87 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1698); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1700 = 8'h88 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1699); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1701 = 8'h89 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1700); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1702 = 8'h8a == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1701); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1703 = 8'h8b == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1702); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1704 = 8'h8c == _GEN_8950 ? $signed(regsA_70_im) : $signed(_GEN_1703); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1705 = 8'h8d == _GEN_8950 ? $signed(regsA_71_im) : $signed(_GEN_1704); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1706 = 8'h8e == _GEN_8950 ? $signed(regsA_72_im) : $signed(_GEN_1705); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1707 = 8'h8f == _GEN_8950 ? $signed(regsA_73_im) : $signed(_GEN_1706); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1708 = 8'h90 == _GEN_8950 ? $signed(regsA_74_im) : $signed(_GEN_1707); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1709 = 8'h91 == _GEN_8950 ? $signed(regsA_75_im) : $signed(_GEN_1708); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1710 = 8'h92 == _GEN_8950 ? $signed(regsA_76_im) : $signed(_GEN_1709); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1711 = 8'h93 == _GEN_8950 ? $signed(regsA_77_im) : $signed(_GEN_1710); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1712 = 8'h94 == _GEN_8950 ? $signed(regsA_78_im) : $signed(_GEN_1711); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1713 = 8'h95 == _GEN_8950 ? $signed(regsA_79_im) : $signed(_GEN_1712); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1714 = 8'h96 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1713); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1715 = 8'h97 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1714); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1716 = 8'h98 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1715); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1717 = 8'h99 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1716); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1718 = 8'h9a == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1717); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1719 = 8'h9b == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1718); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1720 = 8'h9c == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1719); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1721 = 8'h9d == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1720); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1722 = 8'h9e == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1721); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1723 = 8'h9f == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1722); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1724 = 8'ha0 == _GEN_8950 ? $signed(regsA_80_im) : $signed(_GEN_1723); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1725 = 8'ha1 == _GEN_8950 ? $signed(regsA_81_im) : $signed(_GEN_1724); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1726 = 8'ha2 == _GEN_8950 ? $signed(regsA_82_im) : $signed(_GEN_1725); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1727 = 8'ha3 == _GEN_8950 ? $signed(regsA_83_im) : $signed(_GEN_1726); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1728 = 8'ha4 == _GEN_8950 ? $signed(regsA_84_im) : $signed(_GEN_1727); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1729 = 8'ha5 == _GEN_8950 ? $signed(regsA_85_im) : $signed(_GEN_1728); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1730 = 8'ha6 == _GEN_8950 ? $signed(regsA_86_im) : $signed(_GEN_1729); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1731 = 8'ha7 == _GEN_8950 ? $signed(regsA_87_im) : $signed(_GEN_1730); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1732 = 8'ha8 == _GEN_8950 ? $signed(regsA_88_im) : $signed(_GEN_1731); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1733 = 8'ha9 == _GEN_8950 ? $signed(regsA_89_im) : $signed(_GEN_1732); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1734 = 8'haa == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1733); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1735 = 8'hab == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1734); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1736 = 8'hac == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1735); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1737 = 8'had == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1736); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1738 = 8'hae == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1737); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1739 = 8'haf == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1738); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1740 = 8'hb0 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1739); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1741 = 8'hb1 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1740); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1742 = 8'hb2 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1741); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1743 = 8'hb3 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1742); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1744 = 8'hb4 == _GEN_8950 ? $signed(regsA_90_im) : $signed(_GEN_1743); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1745 = 8'hb5 == _GEN_8950 ? $signed(regsA_91_im) : $signed(_GEN_1744); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1746 = 8'hb6 == _GEN_8950 ? $signed(regsA_92_im) : $signed(_GEN_1745); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1747 = 8'hb7 == _GEN_8950 ? $signed(regsA_93_im) : $signed(_GEN_1746); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1748 = 8'hb8 == _GEN_8950 ? $signed(regsA_94_im) : $signed(_GEN_1747); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1749 = 8'hb9 == _GEN_8950 ? $signed(regsA_95_im) : $signed(_GEN_1748); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1750 = 8'hba == _GEN_8950 ? $signed(regsA_96_im) : $signed(_GEN_1749); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1751 = 8'hbb == _GEN_8950 ? $signed(regsA_97_im) : $signed(_GEN_1750); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1752 = 8'hbc == _GEN_8950 ? $signed(regsA_98_im) : $signed(_GEN_1751); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1753 = 8'hbd == _GEN_8950 ? $signed(regsA_99_im) : $signed(_GEN_1752); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1755 = 7'h1 == _T_9 ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1756 = 7'h2 == _T_9 ? $signed(regsA_2_re) : $signed(_GEN_1755); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1757 = 7'h3 == _T_9 ? $signed(regsA_3_re) : $signed(_GEN_1756); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1758 = 7'h4 == _T_9 ? $signed(regsA_4_re) : $signed(_GEN_1757); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1759 = 7'h5 == _T_9 ? $signed(regsA_5_re) : $signed(_GEN_1758); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1760 = 7'h6 == _T_9 ? $signed(regsA_6_re) : $signed(_GEN_1759); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1761 = 7'h7 == _T_9 ? $signed(regsA_7_re) : $signed(_GEN_1760); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1762 = 7'h8 == _T_9 ? $signed(regsA_8_re) : $signed(_GEN_1761); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1763 = 7'h9 == _T_9 ? $signed(regsA_9_re) : $signed(_GEN_1762); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1764 = 7'ha == _T_9 ? $signed(32'sh0) : $signed(_GEN_1763); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1765 = 7'hb == _T_9 ? $signed(32'sh0) : $signed(_GEN_1764); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1766 = 7'hc == _T_9 ? $signed(32'sh0) : $signed(_GEN_1765); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1767 = 7'hd == _T_9 ? $signed(32'sh0) : $signed(_GEN_1766); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1768 = 7'he == _T_9 ? $signed(32'sh0) : $signed(_GEN_1767); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1769 = 7'hf == _T_9 ? $signed(32'sh0) : $signed(_GEN_1768); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1770 = 7'h10 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1769); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1771 = 7'h11 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1770); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1772 = 7'h12 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1771); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1773 = 7'h13 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1772); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1774 = 7'h14 == _T_9 ? $signed(regsA_10_re) : $signed(_GEN_1773); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1775 = 7'h15 == _T_9 ? $signed(regsA_11_re) : $signed(_GEN_1774); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1776 = 7'h16 == _T_9 ? $signed(regsA_12_re) : $signed(_GEN_1775); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1777 = 7'h17 == _T_9 ? $signed(regsA_13_re) : $signed(_GEN_1776); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1778 = 7'h18 == _T_9 ? $signed(regsA_14_re) : $signed(_GEN_1777); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1779 = 7'h19 == _T_9 ? $signed(regsA_15_re) : $signed(_GEN_1778); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1780 = 7'h1a == _T_9 ? $signed(regsA_16_re) : $signed(_GEN_1779); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1781 = 7'h1b == _T_9 ? $signed(regsA_17_re) : $signed(_GEN_1780); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1782 = 7'h1c == _T_9 ? $signed(regsA_18_re) : $signed(_GEN_1781); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1783 = 7'h1d == _T_9 ? $signed(regsA_19_re) : $signed(_GEN_1782); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1784 = 7'h1e == _T_9 ? $signed(32'sh0) : $signed(_GEN_1783); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1785 = 7'h1f == _T_9 ? $signed(32'sh0) : $signed(_GEN_1784); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1786 = 7'h20 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1785); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1787 = 7'h21 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1786); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1788 = 7'h22 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1787); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1789 = 7'h23 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1788); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1790 = 7'h24 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1789); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1791 = 7'h25 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1790); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1792 = 7'h26 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1791); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1793 = 7'h27 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1792); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1794 = 7'h28 == _T_9 ? $signed(regsA_20_re) : $signed(_GEN_1793); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1795 = 7'h29 == _T_9 ? $signed(regsA_21_re) : $signed(_GEN_1794); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1796 = 7'h2a == _T_9 ? $signed(regsA_22_re) : $signed(_GEN_1795); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1797 = 7'h2b == _T_9 ? $signed(regsA_23_re) : $signed(_GEN_1796); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1798 = 7'h2c == _T_9 ? $signed(regsA_24_re) : $signed(_GEN_1797); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1799 = 7'h2d == _T_9 ? $signed(regsA_25_re) : $signed(_GEN_1798); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1800 = 7'h2e == _T_9 ? $signed(regsA_26_re) : $signed(_GEN_1799); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1801 = 7'h2f == _T_9 ? $signed(regsA_27_re) : $signed(_GEN_1800); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1802 = 7'h30 == _T_9 ? $signed(regsA_28_re) : $signed(_GEN_1801); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1803 = 7'h31 == _T_9 ? $signed(regsA_29_re) : $signed(_GEN_1802); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1804 = 7'h32 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1803); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1805 = 7'h33 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1804); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1806 = 7'h34 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1805); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1807 = 7'h35 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1806); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1808 = 7'h36 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1807); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1809 = 7'h37 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1808); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1810 = 7'h38 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1809); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1811 = 7'h39 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1810); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1812 = 7'h3a == _T_9 ? $signed(32'sh0) : $signed(_GEN_1811); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1813 = 7'h3b == _T_9 ? $signed(32'sh0) : $signed(_GEN_1812); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1814 = 7'h3c == _T_9 ? $signed(regsA_30_re) : $signed(_GEN_1813); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1815 = 7'h3d == _T_9 ? $signed(regsA_31_re) : $signed(_GEN_1814); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1816 = 7'h3e == _T_9 ? $signed(regsA_32_re) : $signed(_GEN_1815); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1817 = 7'h3f == _T_9 ? $signed(regsA_33_re) : $signed(_GEN_1816); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1818 = 7'h40 == _T_9 ? $signed(regsA_34_re) : $signed(_GEN_1817); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1819 = 7'h41 == _T_9 ? $signed(regsA_35_re) : $signed(_GEN_1818); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1820 = 7'h42 == _T_9 ? $signed(regsA_36_re) : $signed(_GEN_1819); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1821 = 7'h43 == _T_9 ? $signed(regsA_37_re) : $signed(_GEN_1820); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1822 = 7'h44 == _T_9 ? $signed(regsA_38_re) : $signed(_GEN_1821); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1823 = 7'h45 == _T_9 ? $signed(regsA_39_re) : $signed(_GEN_1822); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1824 = 7'h46 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1823); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1825 = 7'h47 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1824); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1826 = 7'h48 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1825); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1827 = 7'h49 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1826); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1828 = 7'h4a == _T_9 ? $signed(32'sh0) : $signed(_GEN_1827); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1829 = 7'h4b == _T_9 ? $signed(32'sh0) : $signed(_GEN_1828); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1830 = 7'h4c == _T_9 ? $signed(32'sh0) : $signed(_GEN_1829); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1831 = 7'h4d == _T_9 ? $signed(32'sh0) : $signed(_GEN_1830); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1832 = 7'h4e == _T_9 ? $signed(32'sh0) : $signed(_GEN_1831); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1833 = 7'h4f == _T_9 ? $signed(32'sh0) : $signed(_GEN_1832); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1834 = 7'h50 == _T_9 ? $signed(regsA_40_re) : $signed(_GEN_1833); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1835 = 7'h51 == _T_9 ? $signed(regsA_41_re) : $signed(_GEN_1834); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1836 = 7'h52 == _T_9 ? $signed(regsA_42_re) : $signed(_GEN_1835); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1837 = 7'h53 == _T_9 ? $signed(regsA_43_re) : $signed(_GEN_1836); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1838 = 7'h54 == _T_9 ? $signed(regsA_44_re) : $signed(_GEN_1837); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1839 = 7'h55 == _T_9 ? $signed(regsA_45_re) : $signed(_GEN_1838); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1840 = 7'h56 == _T_9 ? $signed(regsA_46_re) : $signed(_GEN_1839); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1841 = 7'h57 == _T_9 ? $signed(regsA_47_re) : $signed(_GEN_1840); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1842 = 7'h58 == _T_9 ? $signed(regsA_48_re) : $signed(_GEN_1841); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1843 = 7'h59 == _T_9 ? $signed(regsA_49_re) : $signed(_GEN_1842); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1844 = 7'h5a == _T_9 ? $signed(32'sh0) : $signed(_GEN_1843); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1845 = 7'h5b == _T_9 ? $signed(32'sh0) : $signed(_GEN_1844); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1846 = 7'h5c == _T_9 ? $signed(32'sh0) : $signed(_GEN_1845); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1847 = 7'h5d == _T_9 ? $signed(32'sh0) : $signed(_GEN_1846); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1848 = 7'h5e == _T_9 ? $signed(32'sh0) : $signed(_GEN_1847); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1849 = 7'h5f == _T_9 ? $signed(32'sh0) : $signed(_GEN_1848); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1850 = 7'h60 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1849); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1851 = 7'h61 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1850); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1852 = 7'h62 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1851); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1853 = 7'h63 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1852); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1854 = 7'h64 == _T_9 ? $signed(regsA_50_re) : $signed(_GEN_1853); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1855 = 7'h65 == _T_9 ? $signed(regsA_51_re) : $signed(_GEN_1854); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1856 = 7'h66 == _T_9 ? $signed(regsA_52_re) : $signed(_GEN_1855); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1857 = 7'h67 == _T_9 ? $signed(regsA_53_re) : $signed(_GEN_1856); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1858 = 7'h68 == _T_9 ? $signed(regsA_54_re) : $signed(_GEN_1857); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1859 = 7'h69 == _T_9 ? $signed(regsA_55_re) : $signed(_GEN_1858); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1860 = 7'h6a == _T_9 ? $signed(regsA_56_re) : $signed(_GEN_1859); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1861 = 7'h6b == _T_9 ? $signed(regsA_57_re) : $signed(_GEN_1860); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1862 = 7'h6c == _T_9 ? $signed(regsA_58_re) : $signed(_GEN_1861); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1863 = 7'h6d == _T_9 ? $signed(regsA_59_re) : $signed(_GEN_1862); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1864 = 7'h6e == _T_9 ? $signed(32'sh0) : $signed(_GEN_1863); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1865 = 7'h6f == _T_9 ? $signed(32'sh0) : $signed(_GEN_1864); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1866 = 7'h70 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1865); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1867 = 7'h71 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1866); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1868 = 7'h72 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1867); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1869 = 7'h73 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1868); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1870 = 7'h74 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1869); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1871 = 7'h75 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1870); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1872 = 7'h76 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1871); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1873 = 7'h77 == _T_9 ? $signed(32'sh0) : $signed(_GEN_1872); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1874 = 7'h78 == _T_9 ? $signed(regsA_60_re) : $signed(_GEN_1873); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1875 = 7'h79 == _T_9 ? $signed(regsA_61_re) : $signed(_GEN_1874); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1876 = 7'h7a == _T_9 ? $signed(regsA_62_re) : $signed(_GEN_1875); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1877 = 7'h7b == _T_9 ? $signed(regsA_63_re) : $signed(_GEN_1876); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1878 = 7'h7c == _T_9 ? $signed(regsA_64_re) : $signed(_GEN_1877); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1879 = 7'h7d == _T_9 ? $signed(regsA_65_re) : $signed(_GEN_1878); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1880 = 7'h7e == _T_9 ? $signed(regsA_66_re) : $signed(_GEN_1879); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1881 = 7'h7f == _T_9 ? $signed(regsA_67_re) : $signed(_GEN_1880); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1882 = 8'h80 == _GEN_8950 ? $signed(regsA_68_re) : $signed(_GEN_1881); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1883 = 8'h81 == _GEN_8950 ? $signed(regsA_69_re) : $signed(_GEN_1882); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1884 = 8'h82 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1883); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1885 = 8'h83 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1884); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1886 = 8'h84 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1885); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1887 = 8'h85 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1886); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1888 = 8'h86 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1887); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1889 = 8'h87 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1888); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1890 = 8'h88 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1889); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1891 = 8'h89 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1890); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1892 = 8'h8a == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1891); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1893 = 8'h8b == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1892); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1894 = 8'h8c == _GEN_8950 ? $signed(regsA_70_re) : $signed(_GEN_1893); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1895 = 8'h8d == _GEN_8950 ? $signed(regsA_71_re) : $signed(_GEN_1894); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1896 = 8'h8e == _GEN_8950 ? $signed(regsA_72_re) : $signed(_GEN_1895); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1897 = 8'h8f == _GEN_8950 ? $signed(regsA_73_re) : $signed(_GEN_1896); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1898 = 8'h90 == _GEN_8950 ? $signed(regsA_74_re) : $signed(_GEN_1897); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1899 = 8'h91 == _GEN_8950 ? $signed(regsA_75_re) : $signed(_GEN_1898); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1900 = 8'h92 == _GEN_8950 ? $signed(regsA_76_re) : $signed(_GEN_1899); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1901 = 8'h93 == _GEN_8950 ? $signed(regsA_77_re) : $signed(_GEN_1900); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1902 = 8'h94 == _GEN_8950 ? $signed(regsA_78_re) : $signed(_GEN_1901); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1903 = 8'h95 == _GEN_8950 ? $signed(regsA_79_re) : $signed(_GEN_1902); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1904 = 8'h96 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1903); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1905 = 8'h97 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1904); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1906 = 8'h98 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1905); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1907 = 8'h99 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1906); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1908 = 8'h9a == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1907); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1909 = 8'h9b == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1908); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1910 = 8'h9c == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1909); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1911 = 8'h9d == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1910); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1912 = 8'h9e == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1911); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1913 = 8'h9f == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1912); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1914 = 8'ha0 == _GEN_8950 ? $signed(regsA_80_re) : $signed(_GEN_1913); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1915 = 8'ha1 == _GEN_8950 ? $signed(regsA_81_re) : $signed(_GEN_1914); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1916 = 8'ha2 == _GEN_8950 ? $signed(regsA_82_re) : $signed(_GEN_1915); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1917 = 8'ha3 == _GEN_8950 ? $signed(regsA_83_re) : $signed(_GEN_1916); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1918 = 8'ha4 == _GEN_8950 ? $signed(regsA_84_re) : $signed(_GEN_1917); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1919 = 8'ha5 == _GEN_8950 ? $signed(regsA_85_re) : $signed(_GEN_1918); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1920 = 8'ha6 == _GEN_8950 ? $signed(regsA_86_re) : $signed(_GEN_1919); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1921 = 8'ha7 == _GEN_8950 ? $signed(regsA_87_re) : $signed(_GEN_1920); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1922 = 8'ha8 == _GEN_8950 ? $signed(regsA_88_re) : $signed(_GEN_1921); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1923 = 8'ha9 == _GEN_8950 ? $signed(regsA_89_re) : $signed(_GEN_1922); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1924 = 8'haa == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1923); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1925 = 8'hab == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1924); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1926 = 8'hac == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1925); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1927 = 8'had == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1926); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1928 = 8'hae == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1927); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1929 = 8'haf == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1928); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1930 = 8'hb0 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1929); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1931 = 8'hb1 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1930); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1932 = 8'hb2 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1931); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1933 = 8'hb3 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_1932); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1934 = 8'hb4 == _GEN_8950 ? $signed(regsA_90_re) : $signed(_GEN_1933); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1935 = 8'hb5 == _GEN_8950 ? $signed(regsA_91_re) : $signed(_GEN_1934); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1936 = 8'hb6 == _GEN_8950 ? $signed(regsA_92_re) : $signed(_GEN_1935); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1937 = 8'hb7 == _GEN_8950 ? $signed(regsA_93_re) : $signed(_GEN_1936); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1938 = 8'hb8 == _GEN_8950 ? $signed(regsA_94_re) : $signed(_GEN_1937); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1939 = 8'hb9 == _GEN_8950 ? $signed(regsA_95_re) : $signed(_GEN_1938); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1940 = 8'hba == _GEN_8950 ? $signed(regsA_96_re) : $signed(_GEN_1939); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1941 = 8'hbb == _GEN_8950 ? $signed(regsA_97_re) : $signed(_GEN_1940); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1942 = 8'hbc == _GEN_8950 ? $signed(regsA_98_re) : $signed(_GEN_1941); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1943 = 8'hbd == _GEN_8950 ? $signed(regsA_99_re) : $signed(_GEN_1942); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [6:0] _T_10 = 2'h3 * 5'h13; // @[Matrix_Mul_V1.scala 148:44]
  wire [6:0] _T_12 = _T_10 + _GEN_8949; // @[Matrix_Mul_V1.scala 148:60]
  wire [31:0] _GEN_1945 = 7'h1 == _T_12 ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1946 = 7'h2 == _T_12 ? $signed(regsA_2_im) : $signed(_GEN_1945); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1947 = 7'h3 == _T_12 ? $signed(regsA_3_im) : $signed(_GEN_1946); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1948 = 7'h4 == _T_12 ? $signed(regsA_4_im) : $signed(_GEN_1947); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1949 = 7'h5 == _T_12 ? $signed(regsA_5_im) : $signed(_GEN_1948); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1950 = 7'h6 == _T_12 ? $signed(regsA_6_im) : $signed(_GEN_1949); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1951 = 7'h7 == _T_12 ? $signed(regsA_7_im) : $signed(_GEN_1950); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1952 = 7'h8 == _T_12 ? $signed(regsA_8_im) : $signed(_GEN_1951); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1953 = 7'h9 == _T_12 ? $signed(regsA_9_im) : $signed(_GEN_1952); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1954 = 7'ha == _T_12 ? $signed(32'sh0) : $signed(_GEN_1953); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1955 = 7'hb == _T_12 ? $signed(32'sh0) : $signed(_GEN_1954); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1956 = 7'hc == _T_12 ? $signed(32'sh0) : $signed(_GEN_1955); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1957 = 7'hd == _T_12 ? $signed(32'sh0) : $signed(_GEN_1956); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1958 = 7'he == _T_12 ? $signed(32'sh0) : $signed(_GEN_1957); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1959 = 7'hf == _T_12 ? $signed(32'sh0) : $signed(_GEN_1958); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1960 = 7'h10 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1959); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1961 = 7'h11 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1960); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1962 = 7'h12 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1961); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1963 = 7'h13 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1962); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1964 = 7'h14 == _T_12 ? $signed(regsA_10_im) : $signed(_GEN_1963); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1965 = 7'h15 == _T_12 ? $signed(regsA_11_im) : $signed(_GEN_1964); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1966 = 7'h16 == _T_12 ? $signed(regsA_12_im) : $signed(_GEN_1965); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1967 = 7'h17 == _T_12 ? $signed(regsA_13_im) : $signed(_GEN_1966); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1968 = 7'h18 == _T_12 ? $signed(regsA_14_im) : $signed(_GEN_1967); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1969 = 7'h19 == _T_12 ? $signed(regsA_15_im) : $signed(_GEN_1968); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1970 = 7'h1a == _T_12 ? $signed(regsA_16_im) : $signed(_GEN_1969); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1971 = 7'h1b == _T_12 ? $signed(regsA_17_im) : $signed(_GEN_1970); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1972 = 7'h1c == _T_12 ? $signed(regsA_18_im) : $signed(_GEN_1971); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1973 = 7'h1d == _T_12 ? $signed(regsA_19_im) : $signed(_GEN_1972); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1974 = 7'h1e == _T_12 ? $signed(32'sh0) : $signed(_GEN_1973); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1975 = 7'h1f == _T_12 ? $signed(32'sh0) : $signed(_GEN_1974); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1976 = 7'h20 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1975); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1977 = 7'h21 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1976); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1978 = 7'h22 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1977); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1979 = 7'h23 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1978); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1980 = 7'h24 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1979); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1981 = 7'h25 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1980); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1982 = 7'h26 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1981); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1983 = 7'h27 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1982); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1984 = 7'h28 == _T_12 ? $signed(regsA_20_im) : $signed(_GEN_1983); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1985 = 7'h29 == _T_12 ? $signed(regsA_21_im) : $signed(_GEN_1984); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1986 = 7'h2a == _T_12 ? $signed(regsA_22_im) : $signed(_GEN_1985); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1987 = 7'h2b == _T_12 ? $signed(regsA_23_im) : $signed(_GEN_1986); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1988 = 7'h2c == _T_12 ? $signed(regsA_24_im) : $signed(_GEN_1987); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1989 = 7'h2d == _T_12 ? $signed(regsA_25_im) : $signed(_GEN_1988); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1990 = 7'h2e == _T_12 ? $signed(regsA_26_im) : $signed(_GEN_1989); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1991 = 7'h2f == _T_12 ? $signed(regsA_27_im) : $signed(_GEN_1990); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1992 = 7'h30 == _T_12 ? $signed(regsA_28_im) : $signed(_GEN_1991); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1993 = 7'h31 == _T_12 ? $signed(regsA_29_im) : $signed(_GEN_1992); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1994 = 7'h32 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1993); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1995 = 7'h33 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1994); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1996 = 7'h34 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1995); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1997 = 7'h35 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1996); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1998 = 7'h36 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1997); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_1999 = 7'h37 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1998); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2000 = 7'h38 == _T_12 ? $signed(32'sh0) : $signed(_GEN_1999); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2001 = 7'h39 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2000); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2002 = 7'h3a == _T_12 ? $signed(32'sh0) : $signed(_GEN_2001); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2003 = 7'h3b == _T_12 ? $signed(32'sh0) : $signed(_GEN_2002); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2004 = 7'h3c == _T_12 ? $signed(regsA_30_im) : $signed(_GEN_2003); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2005 = 7'h3d == _T_12 ? $signed(regsA_31_im) : $signed(_GEN_2004); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2006 = 7'h3e == _T_12 ? $signed(regsA_32_im) : $signed(_GEN_2005); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2007 = 7'h3f == _T_12 ? $signed(regsA_33_im) : $signed(_GEN_2006); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2008 = 7'h40 == _T_12 ? $signed(regsA_34_im) : $signed(_GEN_2007); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2009 = 7'h41 == _T_12 ? $signed(regsA_35_im) : $signed(_GEN_2008); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2010 = 7'h42 == _T_12 ? $signed(regsA_36_im) : $signed(_GEN_2009); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2011 = 7'h43 == _T_12 ? $signed(regsA_37_im) : $signed(_GEN_2010); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2012 = 7'h44 == _T_12 ? $signed(regsA_38_im) : $signed(_GEN_2011); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2013 = 7'h45 == _T_12 ? $signed(regsA_39_im) : $signed(_GEN_2012); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2014 = 7'h46 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2013); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2015 = 7'h47 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2014); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2016 = 7'h48 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2015); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2017 = 7'h49 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2016); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2018 = 7'h4a == _T_12 ? $signed(32'sh0) : $signed(_GEN_2017); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2019 = 7'h4b == _T_12 ? $signed(32'sh0) : $signed(_GEN_2018); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2020 = 7'h4c == _T_12 ? $signed(32'sh0) : $signed(_GEN_2019); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2021 = 7'h4d == _T_12 ? $signed(32'sh0) : $signed(_GEN_2020); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2022 = 7'h4e == _T_12 ? $signed(32'sh0) : $signed(_GEN_2021); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2023 = 7'h4f == _T_12 ? $signed(32'sh0) : $signed(_GEN_2022); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2024 = 7'h50 == _T_12 ? $signed(regsA_40_im) : $signed(_GEN_2023); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2025 = 7'h51 == _T_12 ? $signed(regsA_41_im) : $signed(_GEN_2024); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2026 = 7'h52 == _T_12 ? $signed(regsA_42_im) : $signed(_GEN_2025); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2027 = 7'h53 == _T_12 ? $signed(regsA_43_im) : $signed(_GEN_2026); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2028 = 7'h54 == _T_12 ? $signed(regsA_44_im) : $signed(_GEN_2027); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2029 = 7'h55 == _T_12 ? $signed(regsA_45_im) : $signed(_GEN_2028); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2030 = 7'h56 == _T_12 ? $signed(regsA_46_im) : $signed(_GEN_2029); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2031 = 7'h57 == _T_12 ? $signed(regsA_47_im) : $signed(_GEN_2030); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2032 = 7'h58 == _T_12 ? $signed(regsA_48_im) : $signed(_GEN_2031); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2033 = 7'h59 == _T_12 ? $signed(regsA_49_im) : $signed(_GEN_2032); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2034 = 7'h5a == _T_12 ? $signed(32'sh0) : $signed(_GEN_2033); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2035 = 7'h5b == _T_12 ? $signed(32'sh0) : $signed(_GEN_2034); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2036 = 7'h5c == _T_12 ? $signed(32'sh0) : $signed(_GEN_2035); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2037 = 7'h5d == _T_12 ? $signed(32'sh0) : $signed(_GEN_2036); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2038 = 7'h5e == _T_12 ? $signed(32'sh0) : $signed(_GEN_2037); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2039 = 7'h5f == _T_12 ? $signed(32'sh0) : $signed(_GEN_2038); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2040 = 7'h60 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2039); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2041 = 7'h61 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2040); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2042 = 7'h62 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2041); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2043 = 7'h63 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2042); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2044 = 7'h64 == _T_12 ? $signed(regsA_50_im) : $signed(_GEN_2043); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2045 = 7'h65 == _T_12 ? $signed(regsA_51_im) : $signed(_GEN_2044); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2046 = 7'h66 == _T_12 ? $signed(regsA_52_im) : $signed(_GEN_2045); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2047 = 7'h67 == _T_12 ? $signed(regsA_53_im) : $signed(_GEN_2046); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2048 = 7'h68 == _T_12 ? $signed(regsA_54_im) : $signed(_GEN_2047); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2049 = 7'h69 == _T_12 ? $signed(regsA_55_im) : $signed(_GEN_2048); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2050 = 7'h6a == _T_12 ? $signed(regsA_56_im) : $signed(_GEN_2049); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2051 = 7'h6b == _T_12 ? $signed(regsA_57_im) : $signed(_GEN_2050); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2052 = 7'h6c == _T_12 ? $signed(regsA_58_im) : $signed(_GEN_2051); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2053 = 7'h6d == _T_12 ? $signed(regsA_59_im) : $signed(_GEN_2052); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2054 = 7'h6e == _T_12 ? $signed(32'sh0) : $signed(_GEN_2053); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2055 = 7'h6f == _T_12 ? $signed(32'sh0) : $signed(_GEN_2054); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2056 = 7'h70 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2055); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2057 = 7'h71 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2056); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2058 = 7'h72 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2057); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2059 = 7'h73 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2058); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2060 = 7'h74 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2059); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2061 = 7'h75 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2060); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2062 = 7'h76 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2061); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2063 = 7'h77 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2062); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2064 = 7'h78 == _T_12 ? $signed(regsA_60_im) : $signed(_GEN_2063); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2065 = 7'h79 == _T_12 ? $signed(regsA_61_im) : $signed(_GEN_2064); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2066 = 7'h7a == _T_12 ? $signed(regsA_62_im) : $signed(_GEN_2065); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2067 = 7'h7b == _T_12 ? $signed(regsA_63_im) : $signed(_GEN_2066); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2068 = 7'h7c == _T_12 ? $signed(regsA_64_im) : $signed(_GEN_2067); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2069 = 7'h7d == _T_12 ? $signed(regsA_65_im) : $signed(_GEN_2068); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2070 = 7'h7e == _T_12 ? $signed(regsA_66_im) : $signed(_GEN_2069); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2071 = 7'h7f == _T_12 ? $signed(regsA_67_im) : $signed(_GEN_2070); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [7:0] _GEN_9075 = {{1'd0}, _T_12}; // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2072 = 8'h80 == _GEN_9075 ? $signed(regsA_68_im) : $signed(_GEN_2071); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2073 = 8'h81 == _GEN_9075 ? $signed(regsA_69_im) : $signed(_GEN_2072); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2074 = 8'h82 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2073); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2075 = 8'h83 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2074); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2076 = 8'h84 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2075); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2077 = 8'h85 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2076); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2078 = 8'h86 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2077); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2079 = 8'h87 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2078); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2080 = 8'h88 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2079); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2081 = 8'h89 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2080); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2082 = 8'h8a == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2081); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2083 = 8'h8b == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2082); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2084 = 8'h8c == _GEN_9075 ? $signed(regsA_70_im) : $signed(_GEN_2083); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2085 = 8'h8d == _GEN_9075 ? $signed(regsA_71_im) : $signed(_GEN_2084); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2086 = 8'h8e == _GEN_9075 ? $signed(regsA_72_im) : $signed(_GEN_2085); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2087 = 8'h8f == _GEN_9075 ? $signed(regsA_73_im) : $signed(_GEN_2086); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2088 = 8'h90 == _GEN_9075 ? $signed(regsA_74_im) : $signed(_GEN_2087); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2089 = 8'h91 == _GEN_9075 ? $signed(regsA_75_im) : $signed(_GEN_2088); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2090 = 8'h92 == _GEN_9075 ? $signed(regsA_76_im) : $signed(_GEN_2089); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2091 = 8'h93 == _GEN_9075 ? $signed(regsA_77_im) : $signed(_GEN_2090); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2092 = 8'h94 == _GEN_9075 ? $signed(regsA_78_im) : $signed(_GEN_2091); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2093 = 8'h95 == _GEN_9075 ? $signed(regsA_79_im) : $signed(_GEN_2092); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2094 = 8'h96 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2093); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2095 = 8'h97 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2094); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2096 = 8'h98 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2095); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2097 = 8'h99 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2096); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2098 = 8'h9a == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2097); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2099 = 8'h9b == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2098); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2100 = 8'h9c == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2099); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2101 = 8'h9d == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2100); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2102 = 8'h9e == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2101); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2103 = 8'h9f == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2102); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2104 = 8'ha0 == _GEN_9075 ? $signed(regsA_80_im) : $signed(_GEN_2103); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2105 = 8'ha1 == _GEN_9075 ? $signed(regsA_81_im) : $signed(_GEN_2104); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2106 = 8'ha2 == _GEN_9075 ? $signed(regsA_82_im) : $signed(_GEN_2105); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2107 = 8'ha3 == _GEN_9075 ? $signed(regsA_83_im) : $signed(_GEN_2106); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2108 = 8'ha4 == _GEN_9075 ? $signed(regsA_84_im) : $signed(_GEN_2107); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2109 = 8'ha5 == _GEN_9075 ? $signed(regsA_85_im) : $signed(_GEN_2108); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2110 = 8'ha6 == _GEN_9075 ? $signed(regsA_86_im) : $signed(_GEN_2109); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2111 = 8'ha7 == _GEN_9075 ? $signed(regsA_87_im) : $signed(_GEN_2110); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2112 = 8'ha8 == _GEN_9075 ? $signed(regsA_88_im) : $signed(_GEN_2111); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2113 = 8'ha9 == _GEN_9075 ? $signed(regsA_89_im) : $signed(_GEN_2112); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2114 = 8'haa == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2113); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2115 = 8'hab == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2114); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2116 = 8'hac == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2115); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2117 = 8'had == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2116); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2118 = 8'hae == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2117); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2119 = 8'haf == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2118); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2120 = 8'hb0 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2119); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2121 = 8'hb1 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2120); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2122 = 8'hb2 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2121); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2123 = 8'hb3 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2122); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2124 = 8'hb4 == _GEN_9075 ? $signed(regsA_90_im) : $signed(_GEN_2123); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2125 = 8'hb5 == _GEN_9075 ? $signed(regsA_91_im) : $signed(_GEN_2124); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2126 = 8'hb6 == _GEN_9075 ? $signed(regsA_92_im) : $signed(_GEN_2125); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2127 = 8'hb7 == _GEN_9075 ? $signed(regsA_93_im) : $signed(_GEN_2126); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2128 = 8'hb8 == _GEN_9075 ? $signed(regsA_94_im) : $signed(_GEN_2127); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2129 = 8'hb9 == _GEN_9075 ? $signed(regsA_95_im) : $signed(_GEN_2128); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2130 = 8'hba == _GEN_9075 ? $signed(regsA_96_im) : $signed(_GEN_2129); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2131 = 8'hbb == _GEN_9075 ? $signed(regsA_97_im) : $signed(_GEN_2130); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2132 = 8'hbc == _GEN_9075 ? $signed(regsA_98_im) : $signed(_GEN_2131); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2133 = 8'hbd == _GEN_9075 ? $signed(regsA_99_im) : $signed(_GEN_2132); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2135 = 7'h1 == _T_12 ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2136 = 7'h2 == _T_12 ? $signed(regsA_2_re) : $signed(_GEN_2135); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2137 = 7'h3 == _T_12 ? $signed(regsA_3_re) : $signed(_GEN_2136); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2138 = 7'h4 == _T_12 ? $signed(regsA_4_re) : $signed(_GEN_2137); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2139 = 7'h5 == _T_12 ? $signed(regsA_5_re) : $signed(_GEN_2138); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2140 = 7'h6 == _T_12 ? $signed(regsA_6_re) : $signed(_GEN_2139); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2141 = 7'h7 == _T_12 ? $signed(regsA_7_re) : $signed(_GEN_2140); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2142 = 7'h8 == _T_12 ? $signed(regsA_8_re) : $signed(_GEN_2141); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2143 = 7'h9 == _T_12 ? $signed(regsA_9_re) : $signed(_GEN_2142); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2144 = 7'ha == _T_12 ? $signed(32'sh0) : $signed(_GEN_2143); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2145 = 7'hb == _T_12 ? $signed(32'sh0) : $signed(_GEN_2144); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2146 = 7'hc == _T_12 ? $signed(32'sh0) : $signed(_GEN_2145); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2147 = 7'hd == _T_12 ? $signed(32'sh0) : $signed(_GEN_2146); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2148 = 7'he == _T_12 ? $signed(32'sh0) : $signed(_GEN_2147); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2149 = 7'hf == _T_12 ? $signed(32'sh0) : $signed(_GEN_2148); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2150 = 7'h10 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2149); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2151 = 7'h11 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2150); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2152 = 7'h12 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2151); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2153 = 7'h13 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2152); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2154 = 7'h14 == _T_12 ? $signed(regsA_10_re) : $signed(_GEN_2153); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2155 = 7'h15 == _T_12 ? $signed(regsA_11_re) : $signed(_GEN_2154); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2156 = 7'h16 == _T_12 ? $signed(regsA_12_re) : $signed(_GEN_2155); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2157 = 7'h17 == _T_12 ? $signed(regsA_13_re) : $signed(_GEN_2156); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2158 = 7'h18 == _T_12 ? $signed(regsA_14_re) : $signed(_GEN_2157); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2159 = 7'h19 == _T_12 ? $signed(regsA_15_re) : $signed(_GEN_2158); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2160 = 7'h1a == _T_12 ? $signed(regsA_16_re) : $signed(_GEN_2159); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2161 = 7'h1b == _T_12 ? $signed(regsA_17_re) : $signed(_GEN_2160); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2162 = 7'h1c == _T_12 ? $signed(regsA_18_re) : $signed(_GEN_2161); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2163 = 7'h1d == _T_12 ? $signed(regsA_19_re) : $signed(_GEN_2162); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2164 = 7'h1e == _T_12 ? $signed(32'sh0) : $signed(_GEN_2163); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2165 = 7'h1f == _T_12 ? $signed(32'sh0) : $signed(_GEN_2164); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2166 = 7'h20 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2165); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2167 = 7'h21 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2166); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2168 = 7'h22 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2167); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2169 = 7'h23 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2168); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2170 = 7'h24 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2169); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2171 = 7'h25 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2170); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2172 = 7'h26 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2171); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2173 = 7'h27 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2172); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2174 = 7'h28 == _T_12 ? $signed(regsA_20_re) : $signed(_GEN_2173); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2175 = 7'h29 == _T_12 ? $signed(regsA_21_re) : $signed(_GEN_2174); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2176 = 7'h2a == _T_12 ? $signed(regsA_22_re) : $signed(_GEN_2175); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2177 = 7'h2b == _T_12 ? $signed(regsA_23_re) : $signed(_GEN_2176); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2178 = 7'h2c == _T_12 ? $signed(regsA_24_re) : $signed(_GEN_2177); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2179 = 7'h2d == _T_12 ? $signed(regsA_25_re) : $signed(_GEN_2178); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2180 = 7'h2e == _T_12 ? $signed(regsA_26_re) : $signed(_GEN_2179); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2181 = 7'h2f == _T_12 ? $signed(regsA_27_re) : $signed(_GEN_2180); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2182 = 7'h30 == _T_12 ? $signed(regsA_28_re) : $signed(_GEN_2181); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2183 = 7'h31 == _T_12 ? $signed(regsA_29_re) : $signed(_GEN_2182); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2184 = 7'h32 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2183); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2185 = 7'h33 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2184); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2186 = 7'h34 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2185); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2187 = 7'h35 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2186); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2188 = 7'h36 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2187); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2189 = 7'h37 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2188); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2190 = 7'h38 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2189); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2191 = 7'h39 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2190); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2192 = 7'h3a == _T_12 ? $signed(32'sh0) : $signed(_GEN_2191); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2193 = 7'h3b == _T_12 ? $signed(32'sh0) : $signed(_GEN_2192); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2194 = 7'h3c == _T_12 ? $signed(regsA_30_re) : $signed(_GEN_2193); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2195 = 7'h3d == _T_12 ? $signed(regsA_31_re) : $signed(_GEN_2194); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2196 = 7'h3e == _T_12 ? $signed(regsA_32_re) : $signed(_GEN_2195); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2197 = 7'h3f == _T_12 ? $signed(regsA_33_re) : $signed(_GEN_2196); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2198 = 7'h40 == _T_12 ? $signed(regsA_34_re) : $signed(_GEN_2197); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2199 = 7'h41 == _T_12 ? $signed(regsA_35_re) : $signed(_GEN_2198); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2200 = 7'h42 == _T_12 ? $signed(regsA_36_re) : $signed(_GEN_2199); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2201 = 7'h43 == _T_12 ? $signed(regsA_37_re) : $signed(_GEN_2200); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2202 = 7'h44 == _T_12 ? $signed(regsA_38_re) : $signed(_GEN_2201); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2203 = 7'h45 == _T_12 ? $signed(regsA_39_re) : $signed(_GEN_2202); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2204 = 7'h46 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2203); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2205 = 7'h47 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2204); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2206 = 7'h48 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2205); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2207 = 7'h49 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2206); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2208 = 7'h4a == _T_12 ? $signed(32'sh0) : $signed(_GEN_2207); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2209 = 7'h4b == _T_12 ? $signed(32'sh0) : $signed(_GEN_2208); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2210 = 7'h4c == _T_12 ? $signed(32'sh0) : $signed(_GEN_2209); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2211 = 7'h4d == _T_12 ? $signed(32'sh0) : $signed(_GEN_2210); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2212 = 7'h4e == _T_12 ? $signed(32'sh0) : $signed(_GEN_2211); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2213 = 7'h4f == _T_12 ? $signed(32'sh0) : $signed(_GEN_2212); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2214 = 7'h50 == _T_12 ? $signed(regsA_40_re) : $signed(_GEN_2213); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2215 = 7'h51 == _T_12 ? $signed(regsA_41_re) : $signed(_GEN_2214); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2216 = 7'h52 == _T_12 ? $signed(regsA_42_re) : $signed(_GEN_2215); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2217 = 7'h53 == _T_12 ? $signed(regsA_43_re) : $signed(_GEN_2216); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2218 = 7'h54 == _T_12 ? $signed(regsA_44_re) : $signed(_GEN_2217); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2219 = 7'h55 == _T_12 ? $signed(regsA_45_re) : $signed(_GEN_2218); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2220 = 7'h56 == _T_12 ? $signed(regsA_46_re) : $signed(_GEN_2219); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2221 = 7'h57 == _T_12 ? $signed(regsA_47_re) : $signed(_GEN_2220); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2222 = 7'h58 == _T_12 ? $signed(regsA_48_re) : $signed(_GEN_2221); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2223 = 7'h59 == _T_12 ? $signed(regsA_49_re) : $signed(_GEN_2222); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2224 = 7'h5a == _T_12 ? $signed(32'sh0) : $signed(_GEN_2223); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2225 = 7'h5b == _T_12 ? $signed(32'sh0) : $signed(_GEN_2224); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2226 = 7'h5c == _T_12 ? $signed(32'sh0) : $signed(_GEN_2225); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2227 = 7'h5d == _T_12 ? $signed(32'sh0) : $signed(_GEN_2226); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2228 = 7'h5e == _T_12 ? $signed(32'sh0) : $signed(_GEN_2227); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2229 = 7'h5f == _T_12 ? $signed(32'sh0) : $signed(_GEN_2228); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2230 = 7'h60 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2229); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2231 = 7'h61 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2230); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2232 = 7'h62 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2231); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2233 = 7'h63 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2232); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2234 = 7'h64 == _T_12 ? $signed(regsA_50_re) : $signed(_GEN_2233); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2235 = 7'h65 == _T_12 ? $signed(regsA_51_re) : $signed(_GEN_2234); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2236 = 7'h66 == _T_12 ? $signed(regsA_52_re) : $signed(_GEN_2235); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2237 = 7'h67 == _T_12 ? $signed(regsA_53_re) : $signed(_GEN_2236); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2238 = 7'h68 == _T_12 ? $signed(regsA_54_re) : $signed(_GEN_2237); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2239 = 7'h69 == _T_12 ? $signed(regsA_55_re) : $signed(_GEN_2238); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2240 = 7'h6a == _T_12 ? $signed(regsA_56_re) : $signed(_GEN_2239); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2241 = 7'h6b == _T_12 ? $signed(regsA_57_re) : $signed(_GEN_2240); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2242 = 7'h6c == _T_12 ? $signed(regsA_58_re) : $signed(_GEN_2241); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2243 = 7'h6d == _T_12 ? $signed(regsA_59_re) : $signed(_GEN_2242); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2244 = 7'h6e == _T_12 ? $signed(32'sh0) : $signed(_GEN_2243); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2245 = 7'h6f == _T_12 ? $signed(32'sh0) : $signed(_GEN_2244); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2246 = 7'h70 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2245); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2247 = 7'h71 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2246); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2248 = 7'h72 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2247); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2249 = 7'h73 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2248); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2250 = 7'h74 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2249); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2251 = 7'h75 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2250); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2252 = 7'h76 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2251); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2253 = 7'h77 == _T_12 ? $signed(32'sh0) : $signed(_GEN_2252); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2254 = 7'h78 == _T_12 ? $signed(regsA_60_re) : $signed(_GEN_2253); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2255 = 7'h79 == _T_12 ? $signed(regsA_61_re) : $signed(_GEN_2254); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2256 = 7'h7a == _T_12 ? $signed(regsA_62_re) : $signed(_GEN_2255); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2257 = 7'h7b == _T_12 ? $signed(regsA_63_re) : $signed(_GEN_2256); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2258 = 7'h7c == _T_12 ? $signed(regsA_64_re) : $signed(_GEN_2257); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2259 = 7'h7d == _T_12 ? $signed(regsA_65_re) : $signed(_GEN_2258); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2260 = 7'h7e == _T_12 ? $signed(regsA_66_re) : $signed(_GEN_2259); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2261 = 7'h7f == _T_12 ? $signed(regsA_67_re) : $signed(_GEN_2260); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2262 = 8'h80 == _GEN_9075 ? $signed(regsA_68_re) : $signed(_GEN_2261); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2263 = 8'h81 == _GEN_9075 ? $signed(regsA_69_re) : $signed(_GEN_2262); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2264 = 8'h82 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2263); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2265 = 8'h83 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2264); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2266 = 8'h84 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2265); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2267 = 8'h85 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2266); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2268 = 8'h86 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2267); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2269 = 8'h87 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2268); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2270 = 8'h88 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2269); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2271 = 8'h89 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2270); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2272 = 8'h8a == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2271); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2273 = 8'h8b == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2272); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2274 = 8'h8c == _GEN_9075 ? $signed(regsA_70_re) : $signed(_GEN_2273); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2275 = 8'h8d == _GEN_9075 ? $signed(regsA_71_re) : $signed(_GEN_2274); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2276 = 8'h8e == _GEN_9075 ? $signed(regsA_72_re) : $signed(_GEN_2275); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2277 = 8'h8f == _GEN_9075 ? $signed(regsA_73_re) : $signed(_GEN_2276); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2278 = 8'h90 == _GEN_9075 ? $signed(regsA_74_re) : $signed(_GEN_2277); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2279 = 8'h91 == _GEN_9075 ? $signed(regsA_75_re) : $signed(_GEN_2278); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2280 = 8'h92 == _GEN_9075 ? $signed(regsA_76_re) : $signed(_GEN_2279); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2281 = 8'h93 == _GEN_9075 ? $signed(regsA_77_re) : $signed(_GEN_2280); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2282 = 8'h94 == _GEN_9075 ? $signed(regsA_78_re) : $signed(_GEN_2281); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2283 = 8'h95 == _GEN_9075 ? $signed(regsA_79_re) : $signed(_GEN_2282); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2284 = 8'h96 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2283); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2285 = 8'h97 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2284); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2286 = 8'h98 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2285); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2287 = 8'h99 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2286); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2288 = 8'h9a == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2287); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2289 = 8'h9b == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2288); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2290 = 8'h9c == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2289); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2291 = 8'h9d == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2290); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2292 = 8'h9e == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2291); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2293 = 8'h9f == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2292); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2294 = 8'ha0 == _GEN_9075 ? $signed(regsA_80_re) : $signed(_GEN_2293); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2295 = 8'ha1 == _GEN_9075 ? $signed(regsA_81_re) : $signed(_GEN_2294); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2296 = 8'ha2 == _GEN_9075 ? $signed(regsA_82_re) : $signed(_GEN_2295); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2297 = 8'ha3 == _GEN_9075 ? $signed(regsA_83_re) : $signed(_GEN_2296); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2298 = 8'ha4 == _GEN_9075 ? $signed(regsA_84_re) : $signed(_GEN_2297); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2299 = 8'ha5 == _GEN_9075 ? $signed(regsA_85_re) : $signed(_GEN_2298); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2300 = 8'ha6 == _GEN_9075 ? $signed(regsA_86_re) : $signed(_GEN_2299); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2301 = 8'ha7 == _GEN_9075 ? $signed(regsA_87_re) : $signed(_GEN_2300); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2302 = 8'ha8 == _GEN_9075 ? $signed(regsA_88_re) : $signed(_GEN_2301); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2303 = 8'ha9 == _GEN_9075 ? $signed(regsA_89_re) : $signed(_GEN_2302); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2304 = 8'haa == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2303); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2305 = 8'hab == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2304); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2306 = 8'hac == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2305); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2307 = 8'had == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2306); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2308 = 8'hae == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2307); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2309 = 8'haf == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2308); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2310 = 8'hb0 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2309); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2311 = 8'hb1 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2310); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2312 = 8'hb2 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2311); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2313 = 8'hb3 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_2312); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2314 = 8'hb4 == _GEN_9075 ? $signed(regsA_90_re) : $signed(_GEN_2313); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2315 = 8'hb5 == _GEN_9075 ? $signed(regsA_91_re) : $signed(_GEN_2314); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2316 = 8'hb6 == _GEN_9075 ? $signed(regsA_92_re) : $signed(_GEN_2315); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2317 = 8'hb7 == _GEN_9075 ? $signed(regsA_93_re) : $signed(_GEN_2316); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2318 = 8'hb8 == _GEN_9075 ? $signed(regsA_94_re) : $signed(_GEN_2317); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2319 = 8'hb9 == _GEN_9075 ? $signed(regsA_95_re) : $signed(_GEN_2318); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2320 = 8'hba == _GEN_9075 ? $signed(regsA_96_re) : $signed(_GEN_2319); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2321 = 8'hbb == _GEN_9075 ? $signed(regsA_97_re) : $signed(_GEN_2320); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2322 = 8'hbc == _GEN_9075 ? $signed(regsA_98_re) : $signed(_GEN_2321); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2323 = 8'hbd == _GEN_9075 ? $signed(regsA_99_re) : $signed(_GEN_2322); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [7:0] _T_13 = 3'h4 * 5'h13; // @[Matrix_Mul_V1.scala 148:44]
  wire [7:0] _GEN_9199 = {{2'd0}, input_point}; // @[Matrix_Mul_V1.scala 148:60]
  wire [7:0] _T_15 = _T_13 + _GEN_9199; // @[Matrix_Mul_V1.scala 148:60]
  wire [31:0] _GEN_2325 = 8'h1 == _T_15 ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2326 = 8'h2 == _T_15 ? $signed(regsA_2_im) : $signed(_GEN_2325); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2327 = 8'h3 == _T_15 ? $signed(regsA_3_im) : $signed(_GEN_2326); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2328 = 8'h4 == _T_15 ? $signed(regsA_4_im) : $signed(_GEN_2327); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2329 = 8'h5 == _T_15 ? $signed(regsA_5_im) : $signed(_GEN_2328); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2330 = 8'h6 == _T_15 ? $signed(regsA_6_im) : $signed(_GEN_2329); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2331 = 8'h7 == _T_15 ? $signed(regsA_7_im) : $signed(_GEN_2330); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2332 = 8'h8 == _T_15 ? $signed(regsA_8_im) : $signed(_GEN_2331); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2333 = 8'h9 == _T_15 ? $signed(regsA_9_im) : $signed(_GEN_2332); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2334 = 8'ha == _T_15 ? $signed(32'sh0) : $signed(_GEN_2333); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2335 = 8'hb == _T_15 ? $signed(32'sh0) : $signed(_GEN_2334); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2336 = 8'hc == _T_15 ? $signed(32'sh0) : $signed(_GEN_2335); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2337 = 8'hd == _T_15 ? $signed(32'sh0) : $signed(_GEN_2336); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2338 = 8'he == _T_15 ? $signed(32'sh0) : $signed(_GEN_2337); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2339 = 8'hf == _T_15 ? $signed(32'sh0) : $signed(_GEN_2338); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2340 = 8'h10 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2339); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2341 = 8'h11 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2340); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2342 = 8'h12 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2341); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2343 = 8'h13 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2342); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2344 = 8'h14 == _T_15 ? $signed(regsA_10_im) : $signed(_GEN_2343); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2345 = 8'h15 == _T_15 ? $signed(regsA_11_im) : $signed(_GEN_2344); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2346 = 8'h16 == _T_15 ? $signed(regsA_12_im) : $signed(_GEN_2345); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2347 = 8'h17 == _T_15 ? $signed(regsA_13_im) : $signed(_GEN_2346); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2348 = 8'h18 == _T_15 ? $signed(regsA_14_im) : $signed(_GEN_2347); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2349 = 8'h19 == _T_15 ? $signed(regsA_15_im) : $signed(_GEN_2348); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2350 = 8'h1a == _T_15 ? $signed(regsA_16_im) : $signed(_GEN_2349); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2351 = 8'h1b == _T_15 ? $signed(regsA_17_im) : $signed(_GEN_2350); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2352 = 8'h1c == _T_15 ? $signed(regsA_18_im) : $signed(_GEN_2351); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2353 = 8'h1d == _T_15 ? $signed(regsA_19_im) : $signed(_GEN_2352); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2354 = 8'h1e == _T_15 ? $signed(32'sh0) : $signed(_GEN_2353); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2355 = 8'h1f == _T_15 ? $signed(32'sh0) : $signed(_GEN_2354); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2356 = 8'h20 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2355); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2357 = 8'h21 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2356); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2358 = 8'h22 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2357); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2359 = 8'h23 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2358); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2360 = 8'h24 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2359); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2361 = 8'h25 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2360); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2362 = 8'h26 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2361); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2363 = 8'h27 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2362); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2364 = 8'h28 == _T_15 ? $signed(regsA_20_im) : $signed(_GEN_2363); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2365 = 8'h29 == _T_15 ? $signed(regsA_21_im) : $signed(_GEN_2364); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2366 = 8'h2a == _T_15 ? $signed(regsA_22_im) : $signed(_GEN_2365); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2367 = 8'h2b == _T_15 ? $signed(regsA_23_im) : $signed(_GEN_2366); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2368 = 8'h2c == _T_15 ? $signed(regsA_24_im) : $signed(_GEN_2367); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2369 = 8'h2d == _T_15 ? $signed(regsA_25_im) : $signed(_GEN_2368); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2370 = 8'h2e == _T_15 ? $signed(regsA_26_im) : $signed(_GEN_2369); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2371 = 8'h2f == _T_15 ? $signed(regsA_27_im) : $signed(_GEN_2370); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2372 = 8'h30 == _T_15 ? $signed(regsA_28_im) : $signed(_GEN_2371); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2373 = 8'h31 == _T_15 ? $signed(regsA_29_im) : $signed(_GEN_2372); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2374 = 8'h32 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2373); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2375 = 8'h33 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2374); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2376 = 8'h34 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2375); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2377 = 8'h35 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2376); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2378 = 8'h36 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2377); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2379 = 8'h37 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2378); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2380 = 8'h38 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2379); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2381 = 8'h39 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2380); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2382 = 8'h3a == _T_15 ? $signed(32'sh0) : $signed(_GEN_2381); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2383 = 8'h3b == _T_15 ? $signed(32'sh0) : $signed(_GEN_2382); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2384 = 8'h3c == _T_15 ? $signed(regsA_30_im) : $signed(_GEN_2383); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2385 = 8'h3d == _T_15 ? $signed(regsA_31_im) : $signed(_GEN_2384); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2386 = 8'h3e == _T_15 ? $signed(regsA_32_im) : $signed(_GEN_2385); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2387 = 8'h3f == _T_15 ? $signed(regsA_33_im) : $signed(_GEN_2386); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2388 = 8'h40 == _T_15 ? $signed(regsA_34_im) : $signed(_GEN_2387); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2389 = 8'h41 == _T_15 ? $signed(regsA_35_im) : $signed(_GEN_2388); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2390 = 8'h42 == _T_15 ? $signed(regsA_36_im) : $signed(_GEN_2389); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2391 = 8'h43 == _T_15 ? $signed(regsA_37_im) : $signed(_GEN_2390); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2392 = 8'h44 == _T_15 ? $signed(regsA_38_im) : $signed(_GEN_2391); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2393 = 8'h45 == _T_15 ? $signed(regsA_39_im) : $signed(_GEN_2392); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2394 = 8'h46 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2393); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2395 = 8'h47 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2394); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2396 = 8'h48 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2395); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2397 = 8'h49 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2396); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2398 = 8'h4a == _T_15 ? $signed(32'sh0) : $signed(_GEN_2397); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2399 = 8'h4b == _T_15 ? $signed(32'sh0) : $signed(_GEN_2398); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2400 = 8'h4c == _T_15 ? $signed(32'sh0) : $signed(_GEN_2399); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2401 = 8'h4d == _T_15 ? $signed(32'sh0) : $signed(_GEN_2400); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2402 = 8'h4e == _T_15 ? $signed(32'sh0) : $signed(_GEN_2401); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2403 = 8'h4f == _T_15 ? $signed(32'sh0) : $signed(_GEN_2402); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2404 = 8'h50 == _T_15 ? $signed(regsA_40_im) : $signed(_GEN_2403); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2405 = 8'h51 == _T_15 ? $signed(regsA_41_im) : $signed(_GEN_2404); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2406 = 8'h52 == _T_15 ? $signed(regsA_42_im) : $signed(_GEN_2405); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2407 = 8'h53 == _T_15 ? $signed(regsA_43_im) : $signed(_GEN_2406); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2408 = 8'h54 == _T_15 ? $signed(regsA_44_im) : $signed(_GEN_2407); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2409 = 8'h55 == _T_15 ? $signed(regsA_45_im) : $signed(_GEN_2408); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2410 = 8'h56 == _T_15 ? $signed(regsA_46_im) : $signed(_GEN_2409); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2411 = 8'h57 == _T_15 ? $signed(regsA_47_im) : $signed(_GEN_2410); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2412 = 8'h58 == _T_15 ? $signed(regsA_48_im) : $signed(_GEN_2411); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2413 = 8'h59 == _T_15 ? $signed(regsA_49_im) : $signed(_GEN_2412); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2414 = 8'h5a == _T_15 ? $signed(32'sh0) : $signed(_GEN_2413); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2415 = 8'h5b == _T_15 ? $signed(32'sh0) : $signed(_GEN_2414); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2416 = 8'h5c == _T_15 ? $signed(32'sh0) : $signed(_GEN_2415); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2417 = 8'h5d == _T_15 ? $signed(32'sh0) : $signed(_GEN_2416); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2418 = 8'h5e == _T_15 ? $signed(32'sh0) : $signed(_GEN_2417); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2419 = 8'h5f == _T_15 ? $signed(32'sh0) : $signed(_GEN_2418); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2420 = 8'h60 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2419); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2421 = 8'h61 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2420); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2422 = 8'h62 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2421); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2423 = 8'h63 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2422); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2424 = 8'h64 == _T_15 ? $signed(regsA_50_im) : $signed(_GEN_2423); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2425 = 8'h65 == _T_15 ? $signed(regsA_51_im) : $signed(_GEN_2424); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2426 = 8'h66 == _T_15 ? $signed(regsA_52_im) : $signed(_GEN_2425); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2427 = 8'h67 == _T_15 ? $signed(regsA_53_im) : $signed(_GEN_2426); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2428 = 8'h68 == _T_15 ? $signed(regsA_54_im) : $signed(_GEN_2427); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2429 = 8'h69 == _T_15 ? $signed(regsA_55_im) : $signed(_GEN_2428); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2430 = 8'h6a == _T_15 ? $signed(regsA_56_im) : $signed(_GEN_2429); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2431 = 8'h6b == _T_15 ? $signed(regsA_57_im) : $signed(_GEN_2430); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2432 = 8'h6c == _T_15 ? $signed(regsA_58_im) : $signed(_GEN_2431); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2433 = 8'h6d == _T_15 ? $signed(regsA_59_im) : $signed(_GEN_2432); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2434 = 8'h6e == _T_15 ? $signed(32'sh0) : $signed(_GEN_2433); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2435 = 8'h6f == _T_15 ? $signed(32'sh0) : $signed(_GEN_2434); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2436 = 8'h70 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2435); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2437 = 8'h71 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2436); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2438 = 8'h72 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2437); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2439 = 8'h73 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2438); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2440 = 8'h74 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2439); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2441 = 8'h75 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2440); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2442 = 8'h76 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2441); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2443 = 8'h77 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2442); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2444 = 8'h78 == _T_15 ? $signed(regsA_60_im) : $signed(_GEN_2443); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2445 = 8'h79 == _T_15 ? $signed(regsA_61_im) : $signed(_GEN_2444); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2446 = 8'h7a == _T_15 ? $signed(regsA_62_im) : $signed(_GEN_2445); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2447 = 8'h7b == _T_15 ? $signed(regsA_63_im) : $signed(_GEN_2446); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2448 = 8'h7c == _T_15 ? $signed(regsA_64_im) : $signed(_GEN_2447); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2449 = 8'h7d == _T_15 ? $signed(regsA_65_im) : $signed(_GEN_2448); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2450 = 8'h7e == _T_15 ? $signed(regsA_66_im) : $signed(_GEN_2449); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2451 = 8'h7f == _T_15 ? $signed(regsA_67_im) : $signed(_GEN_2450); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2452 = 8'h80 == _T_15 ? $signed(regsA_68_im) : $signed(_GEN_2451); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2453 = 8'h81 == _T_15 ? $signed(regsA_69_im) : $signed(_GEN_2452); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2454 = 8'h82 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2453); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2455 = 8'h83 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2454); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2456 = 8'h84 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2455); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2457 = 8'h85 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2456); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2458 = 8'h86 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2457); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2459 = 8'h87 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2458); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2460 = 8'h88 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2459); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2461 = 8'h89 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2460); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2462 = 8'h8a == _T_15 ? $signed(32'sh0) : $signed(_GEN_2461); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2463 = 8'h8b == _T_15 ? $signed(32'sh0) : $signed(_GEN_2462); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2464 = 8'h8c == _T_15 ? $signed(regsA_70_im) : $signed(_GEN_2463); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2465 = 8'h8d == _T_15 ? $signed(regsA_71_im) : $signed(_GEN_2464); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2466 = 8'h8e == _T_15 ? $signed(regsA_72_im) : $signed(_GEN_2465); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2467 = 8'h8f == _T_15 ? $signed(regsA_73_im) : $signed(_GEN_2466); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2468 = 8'h90 == _T_15 ? $signed(regsA_74_im) : $signed(_GEN_2467); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2469 = 8'h91 == _T_15 ? $signed(regsA_75_im) : $signed(_GEN_2468); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2470 = 8'h92 == _T_15 ? $signed(regsA_76_im) : $signed(_GEN_2469); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2471 = 8'h93 == _T_15 ? $signed(regsA_77_im) : $signed(_GEN_2470); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2472 = 8'h94 == _T_15 ? $signed(regsA_78_im) : $signed(_GEN_2471); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2473 = 8'h95 == _T_15 ? $signed(regsA_79_im) : $signed(_GEN_2472); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2474 = 8'h96 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2473); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2475 = 8'h97 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2474); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2476 = 8'h98 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2475); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2477 = 8'h99 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2476); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2478 = 8'h9a == _T_15 ? $signed(32'sh0) : $signed(_GEN_2477); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2479 = 8'h9b == _T_15 ? $signed(32'sh0) : $signed(_GEN_2478); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2480 = 8'h9c == _T_15 ? $signed(32'sh0) : $signed(_GEN_2479); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2481 = 8'h9d == _T_15 ? $signed(32'sh0) : $signed(_GEN_2480); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2482 = 8'h9e == _T_15 ? $signed(32'sh0) : $signed(_GEN_2481); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2483 = 8'h9f == _T_15 ? $signed(32'sh0) : $signed(_GEN_2482); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2484 = 8'ha0 == _T_15 ? $signed(regsA_80_im) : $signed(_GEN_2483); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2485 = 8'ha1 == _T_15 ? $signed(regsA_81_im) : $signed(_GEN_2484); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2486 = 8'ha2 == _T_15 ? $signed(regsA_82_im) : $signed(_GEN_2485); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2487 = 8'ha3 == _T_15 ? $signed(regsA_83_im) : $signed(_GEN_2486); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2488 = 8'ha4 == _T_15 ? $signed(regsA_84_im) : $signed(_GEN_2487); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2489 = 8'ha5 == _T_15 ? $signed(regsA_85_im) : $signed(_GEN_2488); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2490 = 8'ha6 == _T_15 ? $signed(regsA_86_im) : $signed(_GEN_2489); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2491 = 8'ha7 == _T_15 ? $signed(regsA_87_im) : $signed(_GEN_2490); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2492 = 8'ha8 == _T_15 ? $signed(regsA_88_im) : $signed(_GEN_2491); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2493 = 8'ha9 == _T_15 ? $signed(regsA_89_im) : $signed(_GEN_2492); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2494 = 8'haa == _T_15 ? $signed(32'sh0) : $signed(_GEN_2493); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2495 = 8'hab == _T_15 ? $signed(32'sh0) : $signed(_GEN_2494); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2496 = 8'hac == _T_15 ? $signed(32'sh0) : $signed(_GEN_2495); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2497 = 8'had == _T_15 ? $signed(32'sh0) : $signed(_GEN_2496); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2498 = 8'hae == _T_15 ? $signed(32'sh0) : $signed(_GEN_2497); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2499 = 8'haf == _T_15 ? $signed(32'sh0) : $signed(_GEN_2498); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2500 = 8'hb0 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2499); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2501 = 8'hb1 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2500); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2502 = 8'hb2 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2501); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2503 = 8'hb3 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2502); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2504 = 8'hb4 == _T_15 ? $signed(regsA_90_im) : $signed(_GEN_2503); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2505 = 8'hb5 == _T_15 ? $signed(regsA_91_im) : $signed(_GEN_2504); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2506 = 8'hb6 == _T_15 ? $signed(regsA_92_im) : $signed(_GEN_2505); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2507 = 8'hb7 == _T_15 ? $signed(regsA_93_im) : $signed(_GEN_2506); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2508 = 8'hb8 == _T_15 ? $signed(regsA_94_im) : $signed(_GEN_2507); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2509 = 8'hb9 == _T_15 ? $signed(regsA_95_im) : $signed(_GEN_2508); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2510 = 8'hba == _T_15 ? $signed(regsA_96_im) : $signed(_GEN_2509); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2511 = 8'hbb == _T_15 ? $signed(regsA_97_im) : $signed(_GEN_2510); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2512 = 8'hbc == _T_15 ? $signed(regsA_98_im) : $signed(_GEN_2511); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2513 = 8'hbd == _T_15 ? $signed(regsA_99_im) : $signed(_GEN_2512); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2515 = 8'h1 == _T_15 ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2516 = 8'h2 == _T_15 ? $signed(regsA_2_re) : $signed(_GEN_2515); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2517 = 8'h3 == _T_15 ? $signed(regsA_3_re) : $signed(_GEN_2516); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2518 = 8'h4 == _T_15 ? $signed(regsA_4_re) : $signed(_GEN_2517); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2519 = 8'h5 == _T_15 ? $signed(regsA_5_re) : $signed(_GEN_2518); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2520 = 8'h6 == _T_15 ? $signed(regsA_6_re) : $signed(_GEN_2519); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2521 = 8'h7 == _T_15 ? $signed(regsA_7_re) : $signed(_GEN_2520); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2522 = 8'h8 == _T_15 ? $signed(regsA_8_re) : $signed(_GEN_2521); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2523 = 8'h9 == _T_15 ? $signed(regsA_9_re) : $signed(_GEN_2522); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2524 = 8'ha == _T_15 ? $signed(32'sh0) : $signed(_GEN_2523); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2525 = 8'hb == _T_15 ? $signed(32'sh0) : $signed(_GEN_2524); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2526 = 8'hc == _T_15 ? $signed(32'sh0) : $signed(_GEN_2525); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2527 = 8'hd == _T_15 ? $signed(32'sh0) : $signed(_GEN_2526); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2528 = 8'he == _T_15 ? $signed(32'sh0) : $signed(_GEN_2527); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2529 = 8'hf == _T_15 ? $signed(32'sh0) : $signed(_GEN_2528); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2530 = 8'h10 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2529); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2531 = 8'h11 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2530); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2532 = 8'h12 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2531); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2533 = 8'h13 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2532); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2534 = 8'h14 == _T_15 ? $signed(regsA_10_re) : $signed(_GEN_2533); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2535 = 8'h15 == _T_15 ? $signed(regsA_11_re) : $signed(_GEN_2534); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2536 = 8'h16 == _T_15 ? $signed(regsA_12_re) : $signed(_GEN_2535); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2537 = 8'h17 == _T_15 ? $signed(regsA_13_re) : $signed(_GEN_2536); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2538 = 8'h18 == _T_15 ? $signed(regsA_14_re) : $signed(_GEN_2537); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2539 = 8'h19 == _T_15 ? $signed(regsA_15_re) : $signed(_GEN_2538); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2540 = 8'h1a == _T_15 ? $signed(regsA_16_re) : $signed(_GEN_2539); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2541 = 8'h1b == _T_15 ? $signed(regsA_17_re) : $signed(_GEN_2540); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2542 = 8'h1c == _T_15 ? $signed(regsA_18_re) : $signed(_GEN_2541); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2543 = 8'h1d == _T_15 ? $signed(regsA_19_re) : $signed(_GEN_2542); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2544 = 8'h1e == _T_15 ? $signed(32'sh0) : $signed(_GEN_2543); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2545 = 8'h1f == _T_15 ? $signed(32'sh0) : $signed(_GEN_2544); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2546 = 8'h20 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2545); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2547 = 8'h21 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2546); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2548 = 8'h22 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2547); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2549 = 8'h23 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2548); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2550 = 8'h24 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2549); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2551 = 8'h25 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2550); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2552 = 8'h26 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2551); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2553 = 8'h27 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2552); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2554 = 8'h28 == _T_15 ? $signed(regsA_20_re) : $signed(_GEN_2553); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2555 = 8'h29 == _T_15 ? $signed(regsA_21_re) : $signed(_GEN_2554); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2556 = 8'h2a == _T_15 ? $signed(regsA_22_re) : $signed(_GEN_2555); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2557 = 8'h2b == _T_15 ? $signed(regsA_23_re) : $signed(_GEN_2556); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2558 = 8'h2c == _T_15 ? $signed(regsA_24_re) : $signed(_GEN_2557); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2559 = 8'h2d == _T_15 ? $signed(regsA_25_re) : $signed(_GEN_2558); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2560 = 8'h2e == _T_15 ? $signed(regsA_26_re) : $signed(_GEN_2559); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2561 = 8'h2f == _T_15 ? $signed(regsA_27_re) : $signed(_GEN_2560); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2562 = 8'h30 == _T_15 ? $signed(regsA_28_re) : $signed(_GEN_2561); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2563 = 8'h31 == _T_15 ? $signed(regsA_29_re) : $signed(_GEN_2562); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2564 = 8'h32 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2563); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2565 = 8'h33 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2564); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2566 = 8'h34 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2565); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2567 = 8'h35 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2566); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2568 = 8'h36 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2567); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2569 = 8'h37 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2568); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2570 = 8'h38 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2569); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2571 = 8'h39 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2570); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2572 = 8'h3a == _T_15 ? $signed(32'sh0) : $signed(_GEN_2571); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2573 = 8'h3b == _T_15 ? $signed(32'sh0) : $signed(_GEN_2572); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2574 = 8'h3c == _T_15 ? $signed(regsA_30_re) : $signed(_GEN_2573); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2575 = 8'h3d == _T_15 ? $signed(regsA_31_re) : $signed(_GEN_2574); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2576 = 8'h3e == _T_15 ? $signed(regsA_32_re) : $signed(_GEN_2575); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2577 = 8'h3f == _T_15 ? $signed(regsA_33_re) : $signed(_GEN_2576); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2578 = 8'h40 == _T_15 ? $signed(regsA_34_re) : $signed(_GEN_2577); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2579 = 8'h41 == _T_15 ? $signed(regsA_35_re) : $signed(_GEN_2578); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2580 = 8'h42 == _T_15 ? $signed(regsA_36_re) : $signed(_GEN_2579); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2581 = 8'h43 == _T_15 ? $signed(regsA_37_re) : $signed(_GEN_2580); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2582 = 8'h44 == _T_15 ? $signed(regsA_38_re) : $signed(_GEN_2581); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2583 = 8'h45 == _T_15 ? $signed(regsA_39_re) : $signed(_GEN_2582); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2584 = 8'h46 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2583); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2585 = 8'h47 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2584); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2586 = 8'h48 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2585); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2587 = 8'h49 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2586); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2588 = 8'h4a == _T_15 ? $signed(32'sh0) : $signed(_GEN_2587); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2589 = 8'h4b == _T_15 ? $signed(32'sh0) : $signed(_GEN_2588); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2590 = 8'h4c == _T_15 ? $signed(32'sh0) : $signed(_GEN_2589); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2591 = 8'h4d == _T_15 ? $signed(32'sh0) : $signed(_GEN_2590); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2592 = 8'h4e == _T_15 ? $signed(32'sh0) : $signed(_GEN_2591); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2593 = 8'h4f == _T_15 ? $signed(32'sh0) : $signed(_GEN_2592); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2594 = 8'h50 == _T_15 ? $signed(regsA_40_re) : $signed(_GEN_2593); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2595 = 8'h51 == _T_15 ? $signed(regsA_41_re) : $signed(_GEN_2594); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2596 = 8'h52 == _T_15 ? $signed(regsA_42_re) : $signed(_GEN_2595); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2597 = 8'h53 == _T_15 ? $signed(regsA_43_re) : $signed(_GEN_2596); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2598 = 8'h54 == _T_15 ? $signed(regsA_44_re) : $signed(_GEN_2597); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2599 = 8'h55 == _T_15 ? $signed(regsA_45_re) : $signed(_GEN_2598); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2600 = 8'h56 == _T_15 ? $signed(regsA_46_re) : $signed(_GEN_2599); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2601 = 8'h57 == _T_15 ? $signed(regsA_47_re) : $signed(_GEN_2600); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2602 = 8'h58 == _T_15 ? $signed(regsA_48_re) : $signed(_GEN_2601); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2603 = 8'h59 == _T_15 ? $signed(regsA_49_re) : $signed(_GEN_2602); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2604 = 8'h5a == _T_15 ? $signed(32'sh0) : $signed(_GEN_2603); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2605 = 8'h5b == _T_15 ? $signed(32'sh0) : $signed(_GEN_2604); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2606 = 8'h5c == _T_15 ? $signed(32'sh0) : $signed(_GEN_2605); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2607 = 8'h5d == _T_15 ? $signed(32'sh0) : $signed(_GEN_2606); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2608 = 8'h5e == _T_15 ? $signed(32'sh0) : $signed(_GEN_2607); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2609 = 8'h5f == _T_15 ? $signed(32'sh0) : $signed(_GEN_2608); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2610 = 8'h60 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2609); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2611 = 8'h61 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2610); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2612 = 8'h62 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2611); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2613 = 8'h63 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2612); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2614 = 8'h64 == _T_15 ? $signed(regsA_50_re) : $signed(_GEN_2613); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2615 = 8'h65 == _T_15 ? $signed(regsA_51_re) : $signed(_GEN_2614); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2616 = 8'h66 == _T_15 ? $signed(regsA_52_re) : $signed(_GEN_2615); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2617 = 8'h67 == _T_15 ? $signed(regsA_53_re) : $signed(_GEN_2616); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2618 = 8'h68 == _T_15 ? $signed(regsA_54_re) : $signed(_GEN_2617); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2619 = 8'h69 == _T_15 ? $signed(regsA_55_re) : $signed(_GEN_2618); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2620 = 8'h6a == _T_15 ? $signed(regsA_56_re) : $signed(_GEN_2619); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2621 = 8'h6b == _T_15 ? $signed(regsA_57_re) : $signed(_GEN_2620); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2622 = 8'h6c == _T_15 ? $signed(regsA_58_re) : $signed(_GEN_2621); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2623 = 8'h6d == _T_15 ? $signed(regsA_59_re) : $signed(_GEN_2622); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2624 = 8'h6e == _T_15 ? $signed(32'sh0) : $signed(_GEN_2623); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2625 = 8'h6f == _T_15 ? $signed(32'sh0) : $signed(_GEN_2624); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2626 = 8'h70 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2625); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2627 = 8'h71 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2626); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2628 = 8'h72 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2627); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2629 = 8'h73 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2628); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2630 = 8'h74 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2629); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2631 = 8'h75 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2630); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2632 = 8'h76 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2631); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2633 = 8'h77 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2632); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2634 = 8'h78 == _T_15 ? $signed(regsA_60_re) : $signed(_GEN_2633); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2635 = 8'h79 == _T_15 ? $signed(regsA_61_re) : $signed(_GEN_2634); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2636 = 8'h7a == _T_15 ? $signed(regsA_62_re) : $signed(_GEN_2635); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2637 = 8'h7b == _T_15 ? $signed(regsA_63_re) : $signed(_GEN_2636); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2638 = 8'h7c == _T_15 ? $signed(regsA_64_re) : $signed(_GEN_2637); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2639 = 8'h7d == _T_15 ? $signed(regsA_65_re) : $signed(_GEN_2638); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2640 = 8'h7e == _T_15 ? $signed(regsA_66_re) : $signed(_GEN_2639); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2641 = 8'h7f == _T_15 ? $signed(regsA_67_re) : $signed(_GEN_2640); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2642 = 8'h80 == _T_15 ? $signed(regsA_68_re) : $signed(_GEN_2641); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2643 = 8'h81 == _T_15 ? $signed(regsA_69_re) : $signed(_GEN_2642); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2644 = 8'h82 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2643); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2645 = 8'h83 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2644); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2646 = 8'h84 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2645); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2647 = 8'h85 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2646); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2648 = 8'h86 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2647); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2649 = 8'h87 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2648); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2650 = 8'h88 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2649); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2651 = 8'h89 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2650); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2652 = 8'h8a == _T_15 ? $signed(32'sh0) : $signed(_GEN_2651); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2653 = 8'h8b == _T_15 ? $signed(32'sh0) : $signed(_GEN_2652); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2654 = 8'h8c == _T_15 ? $signed(regsA_70_re) : $signed(_GEN_2653); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2655 = 8'h8d == _T_15 ? $signed(regsA_71_re) : $signed(_GEN_2654); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2656 = 8'h8e == _T_15 ? $signed(regsA_72_re) : $signed(_GEN_2655); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2657 = 8'h8f == _T_15 ? $signed(regsA_73_re) : $signed(_GEN_2656); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2658 = 8'h90 == _T_15 ? $signed(regsA_74_re) : $signed(_GEN_2657); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2659 = 8'h91 == _T_15 ? $signed(regsA_75_re) : $signed(_GEN_2658); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2660 = 8'h92 == _T_15 ? $signed(regsA_76_re) : $signed(_GEN_2659); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2661 = 8'h93 == _T_15 ? $signed(regsA_77_re) : $signed(_GEN_2660); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2662 = 8'h94 == _T_15 ? $signed(regsA_78_re) : $signed(_GEN_2661); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2663 = 8'h95 == _T_15 ? $signed(regsA_79_re) : $signed(_GEN_2662); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2664 = 8'h96 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2663); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2665 = 8'h97 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2664); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2666 = 8'h98 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2665); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2667 = 8'h99 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2666); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2668 = 8'h9a == _T_15 ? $signed(32'sh0) : $signed(_GEN_2667); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2669 = 8'h9b == _T_15 ? $signed(32'sh0) : $signed(_GEN_2668); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2670 = 8'h9c == _T_15 ? $signed(32'sh0) : $signed(_GEN_2669); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2671 = 8'h9d == _T_15 ? $signed(32'sh0) : $signed(_GEN_2670); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2672 = 8'h9e == _T_15 ? $signed(32'sh0) : $signed(_GEN_2671); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2673 = 8'h9f == _T_15 ? $signed(32'sh0) : $signed(_GEN_2672); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2674 = 8'ha0 == _T_15 ? $signed(regsA_80_re) : $signed(_GEN_2673); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2675 = 8'ha1 == _T_15 ? $signed(regsA_81_re) : $signed(_GEN_2674); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2676 = 8'ha2 == _T_15 ? $signed(regsA_82_re) : $signed(_GEN_2675); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2677 = 8'ha3 == _T_15 ? $signed(regsA_83_re) : $signed(_GEN_2676); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2678 = 8'ha4 == _T_15 ? $signed(regsA_84_re) : $signed(_GEN_2677); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2679 = 8'ha5 == _T_15 ? $signed(regsA_85_re) : $signed(_GEN_2678); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2680 = 8'ha6 == _T_15 ? $signed(regsA_86_re) : $signed(_GEN_2679); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2681 = 8'ha7 == _T_15 ? $signed(regsA_87_re) : $signed(_GEN_2680); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2682 = 8'ha8 == _T_15 ? $signed(regsA_88_re) : $signed(_GEN_2681); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2683 = 8'ha9 == _T_15 ? $signed(regsA_89_re) : $signed(_GEN_2682); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2684 = 8'haa == _T_15 ? $signed(32'sh0) : $signed(_GEN_2683); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2685 = 8'hab == _T_15 ? $signed(32'sh0) : $signed(_GEN_2684); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2686 = 8'hac == _T_15 ? $signed(32'sh0) : $signed(_GEN_2685); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2687 = 8'had == _T_15 ? $signed(32'sh0) : $signed(_GEN_2686); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2688 = 8'hae == _T_15 ? $signed(32'sh0) : $signed(_GEN_2687); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2689 = 8'haf == _T_15 ? $signed(32'sh0) : $signed(_GEN_2688); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2690 = 8'hb0 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2689); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2691 = 8'hb1 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2690); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2692 = 8'hb2 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2691); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2693 = 8'hb3 == _T_15 ? $signed(32'sh0) : $signed(_GEN_2692); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2694 = 8'hb4 == _T_15 ? $signed(regsA_90_re) : $signed(_GEN_2693); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2695 = 8'hb5 == _T_15 ? $signed(regsA_91_re) : $signed(_GEN_2694); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2696 = 8'hb6 == _T_15 ? $signed(regsA_92_re) : $signed(_GEN_2695); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2697 = 8'hb7 == _T_15 ? $signed(regsA_93_re) : $signed(_GEN_2696); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2698 = 8'hb8 == _T_15 ? $signed(regsA_94_re) : $signed(_GEN_2697); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2699 = 8'hb9 == _T_15 ? $signed(regsA_95_re) : $signed(_GEN_2698); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2700 = 8'hba == _T_15 ? $signed(regsA_96_re) : $signed(_GEN_2699); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2701 = 8'hbb == _T_15 ? $signed(regsA_97_re) : $signed(_GEN_2700); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2702 = 8'hbc == _T_15 ? $signed(regsA_98_re) : $signed(_GEN_2701); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2703 = 8'hbd == _T_15 ? $signed(regsA_99_re) : $signed(_GEN_2702); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [7:0] _T_16 = 3'h5 * 5'h13; // @[Matrix_Mul_V1.scala 148:44]
  wire [7:0] _T_18 = _T_16 + _GEN_9199; // @[Matrix_Mul_V1.scala 148:60]
  wire [31:0] _GEN_2705 = 8'h1 == _T_18 ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2706 = 8'h2 == _T_18 ? $signed(regsA_2_im) : $signed(_GEN_2705); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2707 = 8'h3 == _T_18 ? $signed(regsA_3_im) : $signed(_GEN_2706); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2708 = 8'h4 == _T_18 ? $signed(regsA_4_im) : $signed(_GEN_2707); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2709 = 8'h5 == _T_18 ? $signed(regsA_5_im) : $signed(_GEN_2708); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2710 = 8'h6 == _T_18 ? $signed(regsA_6_im) : $signed(_GEN_2709); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2711 = 8'h7 == _T_18 ? $signed(regsA_7_im) : $signed(_GEN_2710); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2712 = 8'h8 == _T_18 ? $signed(regsA_8_im) : $signed(_GEN_2711); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2713 = 8'h9 == _T_18 ? $signed(regsA_9_im) : $signed(_GEN_2712); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2714 = 8'ha == _T_18 ? $signed(32'sh0) : $signed(_GEN_2713); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2715 = 8'hb == _T_18 ? $signed(32'sh0) : $signed(_GEN_2714); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2716 = 8'hc == _T_18 ? $signed(32'sh0) : $signed(_GEN_2715); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2717 = 8'hd == _T_18 ? $signed(32'sh0) : $signed(_GEN_2716); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2718 = 8'he == _T_18 ? $signed(32'sh0) : $signed(_GEN_2717); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2719 = 8'hf == _T_18 ? $signed(32'sh0) : $signed(_GEN_2718); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2720 = 8'h10 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2719); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2721 = 8'h11 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2720); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2722 = 8'h12 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2721); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2723 = 8'h13 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2722); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2724 = 8'h14 == _T_18 ? $signed(regsA_10_im) : $signed(_GEN_2723); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2725 = 8'h15 == _T_18 ? $signed(regsA_11_im) : $signed(_GEN_2724); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2726 = 8'h16 == _T_18 ? $signed(regsA_12_im) : $signed(_GEN_2725); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2727 = 8'h17 == _T_18 ? $signed(regsA_13_im) : $signed(_GEN_2726); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2728 = 8'h18 == _T_18 ? $signed(regsA_14_im) : $signed(_GEN_2727); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2729 = 8'h19 == _T_18 ? $signed(regsA_15_im) : $signed(_GEN_2728); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2730 = 8'h1a == _T_18 ? $signed(regsA_16_im) : $signed(_GEN_2729); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2731 = 8'h1b == _T_18 ? $signed(regsA_17_im) : $signed(_GEN_2730); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2732 = 8'h1c == _T_18 ? $signed(regsA_18_im) : $signed(_GEN_2731); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2733 = 8'h1d == _T_18 ? $signed(regsA_19_im) : $signed(_GEN_2732); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2734 = 8'h1e == _T_18 ? $signed(32'sh0) : $signed(_GEN_2733); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2735 = 8'h1f == _T_18 ? $signed(32'sh0) : $signed(_GEN_2734); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2736 = 8'h20 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2735); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2737 = 8'h21 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2736); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2738 = 8'h22 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2737); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2739 = 8'h23 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2738); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2740 = 8'h24 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2739); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2741 = 8'h25 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2740); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2742 = 8'h26 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2741); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2743 = 8'h27 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2742); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2744 = 8'h28 == _T_18 ? $signed(regsA_20_im) : $signed(_GEN_2743); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2745 = 8'h29 == _T_18 ? $signed(regsA_21_im) : $signed(_GEN_2744); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2746 = 8'h2a == _T_18 ? $signed(regsA_22_im) : $signed(_GEN_2745); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2747 = 8'h2b == _T_18 ? $signed(regsA_23_im) : $signed(_GEN_2746); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2748 = 8'h2c == _T_18 ? $signed(regsA_24_im) : $signed(_GEN_2747); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2749 = 8'h2d == _T_18 ? $signed(regsA_25_im) : $signed(_GEN_2748); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2750 = 8'h2e == _T_18 ? $signed(regsA_26_im) : $signed(_GEN_2749); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2751 = 8'h2f == _T_18 ? $signed(regsA_27_im) : $signed(_GEN_2750); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2752 = 8'h30 == _T_18 ? $signed(regsA_28_im) : $signed(_GEN_2751); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2753 = 8'h31 == _T_18 ? $signed(regsA_29_im) : $signed(_GEN_2752); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2754 = 8'h32 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2753); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2755 = 8'h33 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2754); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2756 = 8'h34 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2755); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2757 = 8'h35 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2756); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2758 = 8'h36 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2757); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2759 = 8'h37 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2758); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2760 = 8'h38 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2759); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2761 = 8'h39 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2760); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2762 = 8'h3a == _T_18 ? $signed(32'sh0) : $signed(_GEN_2761); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2763 = 8'h3b == _T_18 ? $signed(32'sh0) : $signed(_GEN_2762); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2764 = 8'h3c == _T_18 ? $signed(regsA_30_im) : $signed(_GEN_2763); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2765 = 8'h3d == _T_18 ? $signed(regsA_31_im) : $signed(_GEN_2764); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2766 = 8'h3e == _T_18 ? $signed(regsA_32_im) : $signed(_GEN_2765); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2767 = 8'h3f == _T_18 ? $signed(regsA_33_im) : $signed(_GEN_2766); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2768 = 8'h40 == _T_18 ? $signed(regsA_34_im) : $signed(_GEN_2767); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2769 = 8'h41 == _T_18 ? $signed(regsA_35_im) : $signed(_GEN_2768); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2770 = 8'h42 == _T_18 ? $signed(regsA_36_im) : $signed(_GEN_2769); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2771 = 8'h43 == _T_18 ? $signed(regsA_37_im) : $signed(_GEN_2770); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2772 = 8'h44 == _T_18 ? $signed(regsA_38_im) : $signed(_GEN_2771); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2773 = 8'h45 == _T_18 ? $signed(regsA_39_im) : $signed(_GEN_2772); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2774 = 8'h46 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2773); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2775 = 8'h47 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2774); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2776 = 8'h48 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2775); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2777 = 8'h49 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2776); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2778 = 8'h4a == _T_18 ? $signed(32'sh0) : $signed(_GEN_2777); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2779 = 8'h4b == _T_18 ? $signed(32'sh0) : $signed(_GEN_2778); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2780 = 8'h4c == _T_18 ? $signed(32'sh0) : $signed(_GEN_2779); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2781 = 8'h4d == _T_18 ? $signed(32'sh0) : $signed(_GEN_2780); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2782 = 8'h4e == _T_18 ? $signed(32'sh0) : $signed(_GEN_2781); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2783 = 8'h4f == _T_18 ? $signed(32'sh0) : $signed(_GEN_2782); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2784 = 8'h50 == _T_18 ? $signed(regsA_40_im) : $signed(_GEN_2783); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2785 = 8'h51 == _T_18 ? $signed(regsA_41_im) : $signed(_GEN_2784); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2786 = 8'h52 == _T_18 ? $signed(regsA_42_im) : $signed(_GEN_2785); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2787 = 8'h53 == _T_18 ? $signed(regsA_43_im) : $signed(_GEN_2786); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2788 = 8'h54 == _T_18 ? $signed(regsA_44_im) : $signed(_GEN_2787); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2789 = 8'h55 == _T_18 ? $signed(regsA_45_im) : $signed(_GEN_2788); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2790 = 8'h56 == _T_18 ? $signed(regsA_46_im) : $signed(_GEN_2789); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2791 = 8'h57 == _T_18 ? $signed(regsA_47_im) : $signed(_GEN_2790); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2792 = 8'h58 == _T_18 ? $signed(regsA_48_im) : $signed(_GEN_2791); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2793 = 8'h59 == _T_18 ? $signed(regsA_49_im) : $signed(_GEN_2792); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2794 = 8'h5a == _T_18 ? $signed(32'sh0) : $signed(_GEN_2793); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2795 = 8'h5b == _T_18 ? $signed(32'sh0) : $signed(_GEN_2794); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2796 = 8'h5c == _T_18 ? $signed(32'sh0) : $signed(_GEN_2795); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2797 = 8'h5d == _T_18 ? $signed(32'sh0) : $signed(_GEN_2796); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2798 = 8'h5e == _T_18 ? $signed(32'sh0) : $signed(_GEN_2797); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2799 = 8'h5f == _T_18 ? $signed(32'sh0) : $signed(_GEN_2798); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2800 = 8'h60 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2799); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2801 = 8'h61 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2800); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2802 = 8'h62 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2801); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2803 = 8'h63 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2802); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2804 = 8'h64 == _T_18 ? $signed(regsA_50_im) : $signed(_GEN_2803); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2805 = 8'h65 == _T_18 ? $signed(regsA_51_im) : $signed(_GEN_2804); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2806 = 8'h66 == _T_18 ? $signed(regsA_52_im) : $signed(_GEN_2805); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2807 = 8'h67 == _T_18 ? $signed(regsA_53_im) : $signed(_GEN_2806); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2808 = 8'h68 == _T_18 ? $signed(regsA_54_im) : $signed(_GEN_2807); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2809 = 8'h69 == _T_18 ? $signed(regsA_55_im) : $signed(_GEN_2808); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2810 = 8'h6a == _T_18 ? $signed(regsA_56_im) : $signed(_GEN_2809); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2811 = 8'h6b == _T_18 ? $signed(regsA_57_im) : $signed(_GEN_2810); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2812 = 8'h6c == _T_18 ? $signed(regsA_58_im) : $signed(_GEN_2811); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2813 = 8'h6d == _T_18 ? $signed(regsA_59_im) : $signed(_GEN_2812); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2814 = 8'h6e == _T_18 ? $signed(32'sh0) : $signed(_GEN_2813); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2815 = 8'h6f == _T_18 ? $signed(32'sh0) : $signed(_GEN_2814); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2816 = 8'h70 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2815); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2817 = 8'h71 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2816); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2818 = 8'h72 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2817); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2819 = 8'h73 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2818); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2820 = 8'h74 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2819); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2821 = 8'h75 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2820); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2822 = 8'h76 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2821); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2823 = 8'h77 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2822); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2824 = 8'h78 == _T_18 ? $signed(regsA_60_im) : $signed(_GEN_2823); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2825 = 8'h79 == _T_18 ? $signed(regsA_61_im) : $signed(_GEN_2824); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2826 = 8'h7a == _T_18 ? $signed(regsA_62_im) : $signed(_GEN_2825); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2827 = 8'h7b == _T_18 ? $signed(regsA_63_im) : $signed(_GEN_2826); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2828 = 8'h7c == _T_18 ? $signed(regsA_64_im) : $signed(_GEN_2827); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2829 = 8'h7d == _T_18 ? $signed(regsA_65_im) : $signed(_GEN_2828); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2830 = 8'h7e == _T_18 ? $signed(regsA_66_im) : $signed(_GEN_2829); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2831 = 8'h7f == _T_18 ? $signed(regsA_67_im) : $signed(_GEN_2830); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2832 = 8'h80 == _T_18 ? $signed(regsA_68_im) : $signed(_GEN_2831); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2833 = 8'h81 == _T_18 ? $signed(regsA_69_im) : $signed(_GEN_2832); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2834 = 8'h82 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2833); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2835 = 8'h83 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2834); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2836 = 8'h84 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2835); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2837 = 8'h85 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2836); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2838 = 8'h86 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2837); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2839 = 8'h87 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2838); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2840 = 8'h88 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2839); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2841 = 8'h89 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2840); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2842 = 8'h8a == _T_18 ? $signed(32'sh0) : $signed(_GEN_2841); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2843 = 8'h8b == _T_18 ? $signed(32'sh0) : $signed(_GEN_2842); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2844 = 8'h8c == _T_18 ? $signed(regsA_70_im) : $signed(_GEN_2843); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2845 = 8'h8d == _T_18 ? $signed(regsA_71_im) : $signed(_GEN_2844); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2846 = 8'h8e == _T_18 ? $signed(regsA_72_im) : $signed(_GEN_2845); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2847 = 8'h8f == _T_18 ? $signed(regsA_73_im) : $signed(_GEN_2846); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2848 = 8'h90 == _T_18 ? $signed(regsA_74_im) : $signed(_GEN_2847); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2849 = 8'h91 == _T_18 ? $signed(regsA_75_im) : $signed(_GEN_2848); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2850 = 8'h92 == _T_18 ? $signed(regsA_76_im) : $signed(_GEN_2849); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2851 = 8'h93 == _T_18 ? $signed(regsA_77_im) : $signed(_GEN_2850); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2852 = 8'h94 == _T_18 ? $signed(regsA_78_im) : $signed(_GEN_2851); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2853 = 8'h95 == _T_18 ? $signed(regsA_79_im) : $signed(_GEN_2852); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2854 = 8'h96 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2853); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2855 = 8'h97 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2854); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2856 = 8'h98 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2855); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2857 = 8'h99 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2856); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2858 = 8'h9a == _T_18 ? $signed(32'sh0) : $signed(_GEN_2857); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2859 = 8'h9b == _T_18 ? $signed(32'sh0) : $signed(_GEN_2858); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2860 = 8'h9c == _T_18 ? $signed(32'sh0) : $signed(_GEN_2859); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2861 = 8'h9d == _T_18 ? $signed(32'sh0) : $signed(_GEN_2860); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2862 = 8'h9e == _T_18 ? $signed(32'sh0) : $signed(_GEN_2861); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2863 = 8'h9f == _T_18 ? $signed(32'sh0) : $signed(_GEN_2862); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2864 = 8'ha0 == _T_18 ? $signed(regsA_80_im) : $signed(_GEN_2863); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2865 = 8'ha1 == _T_18 ? $signed(regsA_81_im) : $signed(_GEN_2864); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2866 = 8'ha2 == _T_18 ? $signed(regsA_82_im) : $signed(_GEN_2865); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2867 = 8'ha3 == _T_18 ? $signed(regsA_83_im) : $signed(_GEN_2866); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2868 = 8'ha4 == _T_18 ? $signed(regsA_84_im) : $signed(_GEN_2867); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2869 = 8'ha5 == _T_18 ? $signed(regsA_85_im) : $signed(_GEN_2868); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2870 = 8'ha6 == _T_18 ? $signed(regsA_86_im) : $signed(_GEN_2869); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2871 = 8'ha7 == _T_18 ? $signed(regsA_87_im) : $signed(_GEN_2870); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2872 = 8'ha8 == _T_18 ? $signed(regsA_88_im) : $signed(_GEN_2871); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2873 = 8'ha9 == _T_18 ? $signed(regsA_89_im) : $signed(_GEN_2872); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2874 = 8'haa == _T_18 ? $signed(32'sh0) : $signed(_GEN_2873); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2875 = 8'hab == _T_18 ? $signed(32'sh0) : $signed(_GEN_2874); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2876 = 8'hac == _T_18 ? $signed(32'sh0) : $signed(_GEN_2875); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2877 = 8'had == _T_18 ? $signed(32'sh0) : $signed(_GEN_2876); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2878 = 8'hae == _T_18 ? $signed(32'sh0) : $signed(_GEN_2877); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2879 = 8'haf == _T_18 ? $signed(32'sh0) : $signed(_GEN_2878); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2880 = 8'hb0 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2879); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2881 = 8'hb1 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2880); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2882 = 8'hb2 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2881); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2883 = 8'hb3 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2882); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2884 = 8'hb4 == _T_18 ? $signed(regsA_90_im) : $signed(_GEN_2883); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2885 = 8'hb5 == _T_18 ? $signed(regsA_91_im) : $signed(_GEN_2884); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2886 = 8'hb6 == _T_18 ? $signed(regsA_92_im) : $signed(_GEN_2885); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2887 = 8'hb7 == _T_18 ? $signed(regsA_93_im) : $signed(_GEN_2886); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2888 = 8'hb8 == _T_18 ? $signed(regsA_94_im) : $signed(_GEN_2887); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2889 = 8'hb9 == _T_18 ? $signed(regsA_95_im) : $signed(_GEN_2888); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2890 = 8'hba == _T_18 ? $signed(regsA_96_im) : $signed(_GEN_2889); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2891 = 8'hbb == _T_18 ? $signed(regsA_97_im) : $signed(_GEN_2890); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2892 = 8'hbc == _T_18 ? $signed(regsA_98_im) : $signed(_GEN_2891); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2893 = 8'hbd == _T_18 ? $signed(regsA_99_im) : $signed(_GEN_2892); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2895 = 8'h1 == _T_18 ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2896 = 8'h2 == _T_18 ? $signed(regsA_2_re) : $signed(_GEN_2895); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2897 = 8'h3 == _T_18 ? $signed(regsA_3_re) : $signed(_GEN_2896); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2898 = 8'h4 == _T_18 ? $signed(regsA_4_re) : $signed(_GEN_2897); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2899 = 8'h5 == _T_18 ? $signed(regsA_5_re) : $signed(_GEN_2898); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2900 = 8'h6 == _T_18 ? $signed(regsA_6_re) : $signed(_GEN_2899); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2901 = 8'h7 == _T_18 ? $signed(regsA_7_re) : $signed(_GEN_2900); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2902 = 8'h8 == _T_18 ? $signed(regsA_8_re) : $signed(_GEN_2901); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2903 = 8'h9 == _T_18 ? $signed(regsA_9_re) : $signed(_GEN_2902); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2904 = 8'ha == _T_18 ? $signed(32'sh0) : $signed(_GEN_2903); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2905 = 8'hb == _T_18 ? $signed(32'sh0) : $signed(_GEN_2904); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2906 = 8'hc == _T_18 ? $signed(32'sh0) : $signed(_GEN_2905); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2907 = 8'hd == _T_18 ? $signed(32'sh0) : $signed(_GEN_2906); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2908 = 8'he == _T_18 ? $signed(32'sh0) : $signed(_GEN_2907); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2909 = 8'hf == _T_18 ? $signed(32'sh0) : $signed(_GEN_2908); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2910 = 8'h10 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2909); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2911 = 8'h11 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2910); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2912 = 8'h12 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2911); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2913 = 8'h13 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2912); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2914 = 8'h14 == _T_18 ? $signed(regsA_10_re) : $signed(_GEN_2913); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2915 = 8'h15 == _T_18 ? $signed(regsA_11_re) : $signed(_GEN_2914); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2916 = 8'h16 == _T_18 ? $signed(regsA_12_re) : $signed(_GEN_2915); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2917 = 8'h17 == _T_18 ? $signed(regsA_13_re) : $signed(_GEN_2916); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2918 = 8'h18 == _T_18 ? $signed(regsA_14_re) : $signed(_GEN_2917); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2919 = 8'h19 == _T_18 ? $signed(regsA_15_re) : $signed(_GEN_2918); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2920 = 8'h1a == _T_18 ? $signed(regsA_16_re) : $signed(_GEN_2919); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2921 = 8'h1b == _T_18 ? $signed(regsA_17_re) : $signed(_GEN_2920); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2922 = 8'h1c == _T_18 ? $signed(regsA_18_re) : $signed(_GEN_2921); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2923 = 8'h1d == _T_18 ? $signed(regsA_19_re) : $signed(_GEN_2922); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2924 = 8'h1e == _T_18 ? $signed(32'sh0) : $signed(_GEN_2923); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2925 = 8'h1f == _T_18 ? $signed(32'sh0) : $signed(_GEN_2924); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2926 = 8'h20 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2925); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2927 = 8'h21 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2926); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2928 = 8'h22 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2927); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2929 = 8'h23 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2928); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2930 = 8'h24 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2929); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2931 = 8'h25 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2930); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2932 = 8'h26 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2931); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2933 = 8'h27 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2932); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2934 = 8'h28 == _T_18 ? $signed(regsA_20_re) : $signed(_GEN_2933); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2935 = 8'h29 == _T_18 ? $signed(regsA_21_re) : $signed(_GEN_2934); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2936 = 8'h2a == _T_18 ? $signed(regsA_22_re) : $signed(_GEN_2935); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2937 = 8'h2b == _T_18 ? $signed(regsA_23_re) : $signed(_GEN_2936); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2938 = 8'h2c == _T_18 ? $signed(regsA_24_re) : $signed(_GEN_2937); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2939 = 8'h2d == _T_18 ? $signed(regsA_25_re) : $signed(_GEN_2938); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2940 = 8'h2e == _T_18 ? $signed(regsA_26_re) : $signed(_GEN_2939); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2941 = 8'h2f == _T_18 ? $signed(regsA_27_re) : $signed(_GEN_2940); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2942 = 8'h30 == _T_18 ? $signed(regsA_28_re) : $signed(_GEN_2941); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2943 = 8'h31 == _T_18 ? $signed(regsA_29_re) : $signed(_GEN_2942); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2944 = 8'h32 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2943); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2945 = 8'h33 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2944); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2946 = 8'h34 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2945); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2947 = 8'h35 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2946); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2948 = 8'h36 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2947); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2949 = 8'h37 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2948); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2950 = 8'h38 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2949); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2951 = 8'h39 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2950); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2952 = 8'h3a == _T_18 ? $signed(32'sh0) : $signed(_GEN_2951); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2953 = 8'h3b == _T_18 ? $signed(32'sh0) : $signed(_GEN_2952); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2954 = 8'h3c == _T_18 ? $signed(regsA_30_re) : $signed(_GEN_2953); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2955 = 8'h3d == _T_18 ? $signed(regsA_31_re) : $signed(_GEN_2954); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2956 = 8'h3e == _T_18 ? $signed(regsA_32_re) : $signed(_GEN_2955); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2957 = 8'h3f == _T_18 ? $signed(regsA_33_re) : $signed(_GEN_2956); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2958 = 8'h40 == _T_18 ? $signed(regsA_34_re) : $signed(_GEN_2957); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2959 = 8'h41 == _T_18 ? $signed(regsA_35_re) : $signed(_GEN_2958); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2960 = 8'h42 == _T_18 ? $signed(regsA_36_re) : $signed(_GEN_2959); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2961 = 8'h43 == _T_18 ? $signed(regsA_37_re) : $signed(_GEN_2960); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2962 = 8'h44 == _T_18 ? $signed(regsA_38_re) : $signed(_GEN_2961); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2963 = 8'h45 == _T_18 ? $signed(regsA_39_re) : $signed(_GEN_2962); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2964 = 8'h46 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2963); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2965 = 8'h47 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2964); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2966 = 8'h48 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2965); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2967 = 8'h49 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2966); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2968 = 8'h4a == _T_18 ? $signed(32'sh0) : $signed(_GEN_2967); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2969 = 8'h4b == _T_18 ? $signed(32'sh0) : $signed(_GEN_2968); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2970 = 8'h4c == _T_18 ? $signed(32'sh0) : $signed(_GEN_2969); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2971 = 8'h4d == _T_18 ? $signed(32'sh0) : $signed(_GEN_2970); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2972 = 8'h4e == _T_18 ? $signed(32'sh0) : $signed(_GEN_2971); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2973 = 8'h4f == _T_18 ? $signed(32'sh0) : $signed(_GEN_2972); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2974 = 8'h50 == _T_18 ? $signed(regsA_40_re) : $signed(_GEN_2973); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2975 = 8'h51 == _T_18 ? $signed(regsA_41_re) : $signed(_GEN_2974); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2976 = 8'h52 == _T_18 ? $signed(regsA_42_re) : $signed(_GEN_2975); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2977 = 8'h53 == _T_18 ? $signed(regsA_43_re) : $signed(_GEN_2976); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2978 = 8'h54 == _T_18 ? $signed(regsA_44_re) : $signed(_GEN_2977); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2979 = 8'h55 == _T_18 ? $signed(regsA_45_re) : $signed(_GEN_2978); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2980 = 8'h56 == _T_18 ? $signed(regsA_46_re) : $signed(_GEN_2979); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2981 = 8'h57 == _T_18 ? $signed(regsA_47_re) : $signed(_GEN_2980); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2982 = 8'h58 == _T_18 ? $signed(regsA_48_re) : $signed(_GEN_2981); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2983 = 8'h59 == _T_18 ? $signed(regsA_49_re) : $signed(_GEN_2982); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2984 = 8'h5a == _T_18 ? $signed(32'sh0) : $signed(_GEN_2983); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2985 = 8'h5b == _T_18 ? $signed(32'sh0) : $signed(_GEN_2984); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2986 = 8'h5c == _T_18 ? $signed(32'sh0) : $signed(_GEN_2985); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2987 = 8'h5d == _T_18 ? $signed(32'sh0) : $signed(_GEN_2986); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2988 = 8'h5e == _T_18 ? $signed(32'sh0) : $signed(_GEN_2987); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2989 = 8'h5f == _T_18 ? $signed(32'sh0) : $signed(_GEN_2988); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2990 = 8'h60 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2989); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2991 = 8'h61 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2990); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2992 = 8'h62 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2991); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2993 = 8'h63 == _T_18 ? $signed(32'sh0) : $signed(_GEN_2992); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2994 = 8'h64 == _T_18 ? $signed(regsA_50_re) : $signed(_GEN_2993); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2995 = 8'h65 == _T_18 ? $signed(regsA_51_re) : $signed(_GEN_2994); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2996 = 8'h66 == _T_18 ? $signed(regsA_52_re) : $signed(_GEN_2995); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2997 = 8'h67 == _T_18 ? $signed(regsA_53_re) : $signed(_GEN_2996); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2998 = 8'h68 == _T_18 ? $signed(regsA_54_re) : $signed(_GEN_2997); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_2999 = 8'h69 == _T_18 ? $signed(regsA_55_re) : $signed(_GEN_2998); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3000 = 8'h6a == _T_18 ? $signed(regsA_56_re) : $signed(_GEN_2999); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3001 = 8'h6b == _T_18 ? $signed(regsA_57_re) : $signed(_GEN_3000); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3002 = 8'h6c == _T_18 ? $signed(regsA_58_re) : $signed(_GEN_3001); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3003 = 8'h6d == _T_18 ? $signed(regsA_59_re) : $signed(_GEN_3002); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3004 = 8'h6e == _T_18 ? $signed(32'sh0) : $signed(_GEN_3003); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3005 = 8'h6f == _T_18 ? $signed(32'sh0) : $signed(_GEN_3004); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3006 = 8'h70 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3005); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3007 = 8'h71 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3006); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3008 = 8'h72 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3007); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3009 = 8'h73 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3008); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3010 = 8'h74 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3009); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3011 = 8'h75 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3010); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3012 = 8'h76 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3011); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3013 = 8'h77 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3012); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3014 = 8'h78 == _T_18 ? $signed(regsA_60_re) : $signed(_GEN_3013); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3015 = 8'h79 == _T_18 ? $signed(regsA_61_re) : $signed(_GEN_3014); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3016 = 8'h7a == _T_18 ? $signed(regsA_62_re) : $signed(_GEN_3015); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3017 = 8'h7b == _T_18 ? $signed(regsA_63_re) : $signed(_GEN_3016); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3018 = 8'h7c == _T_18 ? $signed(regsA_64_re) : $signed(_GEN_3017); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3019 = 8'h7d == _T_18 ? $signed(regsA_65_re) : $signed(_GEN_3018); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3020 = 8'h7e == _T_18 ? $signed(regsA_66_re) : $signed(_GEN_3019); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3021 = 8'h7f == _T_18 ? $signed(regsA_67_re) : $signed(_GEN_3020); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3022 = 8'h80 == _T_18 ? $signed(regsA_68_re) : $signed(_GEN_3021); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3023 = 8'h81 == _T_18 ? $signed(regsA_69_re) : $signed(_GEN_3022); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3024 = 8'h82 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3023); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3025 = 8'h83 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3024); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3026 = 8'h84 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3025); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3027 = 8'h85 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3026); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3028 = 8'h86 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3027); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3029 = 8'h87 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3028); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3030 = 8'h88 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3029); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3031 = 8'h89 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3030); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3032 = 8'h8a == _T_18 ? $signed(32'sh0) : $signed(_GEN_3031); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3033 = 8'h8b == _T_18 ? $signed(32'sh0) : $signed(_GEN_3032); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3034 = 8'h8c == _T_18 ? $signed(regsA_70_re) : $signed(_GEN_3033); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3035 = 8'h8d == _T_18 ? $signed(regsA_71_re) : $signed(_GEN_3034); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3036 = 8'h8e == _T_18 ? $signed(regsA_72_re) : $signed(_GEN_3035); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3037 = 8'h8f == _T_18 ? $signed(regsA_73_re) : $signed(_GEN_3036); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3038 = 8'h90 == _T_18 ? $signed(regsA_74_re) : $signed(_GEN_3037); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3039 = 8'h91 == _T_18 ? $signed(regsA_75_re) : $signed(_GEN_3038); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3040 = 8'h92 == _T_18 ? $signed(regsA_76_re) : $signed(_GEN_3039); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3041 = 8'h93 == _T_18 ? $signed(regsA_77_re) : $signed(_GEN_3040); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3042 = 8'h94 == _T_18 ? $signed(regsA_78_re) : $signed(_GEN_3041); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3043 = 8'h95 == _T_18 ? $signed(regsA_79_re) : $signed(_GEN_3042); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3044 = 8'h96 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3043); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3045 = 8'h97 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3044); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3046 = 8'h98 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3045); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3047 = 8'h99 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3046); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3048 = 8'h9a == _T_18 ? $signed(32'sh0) : $signed(_GEN_3047); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3049 = 8'h9b == _T_18 ? $signed(32'sh0) : $signed(_GEN_3048); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3050 = 8'h9c == _T_18 ? $signed(32'sh0) : $signed(_GEN_3049); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3051 = 8'h9d == _T_18 ? $signed(32'sh0) : $signed(_GEN_3050); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3052 = 8'h9e == _T_18 ? $signed(32'sh0) : $signed(_GEN_3051); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3053 = 8'h9f == _T_18 ? $signed(32'sh0) : $signed(_GEN_3052); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3054 = 8'ha0 == _T_18 ? $signed(regsA_80_re) : $signed(_GEN_3053); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3055 = 8'ha1 == _T_18 ? $signed(regsA_81_re) : $signed(_GEN_3054); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3056 = 8'ha2 == _T_18 ? $signed(regsA_82_re) : $signed(_GEN_3055); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3057 = 8'ha3 == _T_18 ? $signed(regsA_83_re) : $signed(_GEN_3056); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3058 = 8'ha4 == _T_18 ? $signed(regsA_84_re) : $signed(_GEN_3057); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3059 = 8'ha5 == _T_18 ? $signed(regsA_85_re) : $signed(_GEN_3058); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3060 = 8'ha6 == _T_18 ? $signed(regsA_86_re) : $signed(_GEN_3059); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3061 = 8'ha7 == _T_18 ? $signed(regsA_87_re) : $signed(_GEN_3060); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3062 = 8'ha8 == _T_18 ? $signed(regsA_88_re) : $signed(_GEN_3061); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3063 = 8'ha9 == _T_18 ? $signed(regsA_89_re) : $signed(_GEN_3062); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3064 = 8'haa == _T_18 ? $signed(32'sh0) : $signed(_GEN_3063); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3065 = 8'hab == _T_18 ? $signed(32'sh0) : $signed(_GEN_3064); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3066 = 8'hac == _T_18 ? $signed(32'sh0) : $signed(_GEN_3065); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3067 = 8'had == _T_18 ? $signed(32'sh0) : $signed(_GEN_3066); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3068 = 8'hae == _T_18 ? $signed(32'sh0) : $signed(_GEN_3067); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3069 = 8'haf == _T_18 ? $signed(32'sh0) : $signed(_GEN_3068); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3070 = 8'hb0 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3069); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3071 = 8'hb1 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3070); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3072 = 8'hb2 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3071); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3073 = 8'hb3 == _T_18 ? $signed(32'sh0) : $signed(_GEN_3072); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3074 = 8'hb4 == _T_18 ? $signed(regsA_90_re) : $signed(_GEN_3073); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3075 = 8'hb5 == _T_18 ? $signed(regsA_91_re) : $signed(_GEN_3074); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3076 = 8'hb6 == _T_18 ? $signed(regsA_92_re) : $signed(_GEN_3075); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3077 = 8'hb7 == _T_18 ? $signed(regsA_93_re) : $signed(_GEN_3076); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3078 = 8'hb8 == _T_18 ? $signed(regsA_94_re) : $signed(_GEN_3077); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3079 = 8'hb9 == _T_18 ? $signed(regsA_95_re) : $signed(_GEN_3078); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3080 = 8'hba == _T_18 ? $signed(regsA_96_re) : $signed(_GEN_3079); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3081 = 8'hbb == _T_18 ? $signed(regsA_97_re) : $signed(_GEN_3080); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3082 = 8'hbc == _T_18 ? $signed(regsA_98_re) : $signed(_GEN_3081); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3083 = 8'hbd == _T_18 ? $signed(regsA_99_re) : $signed(_GEN_3082); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [7:0] _T_19 = 3'h6 * 5'h13; // @[Matrix_Mul_V1.scala 148:44]
  wire [7:0] _T_21 = _T_19 + _GEN_9199; // @[Matrix_Mul_V1.scala 148:60]
  wire [31:0] _GEN_3085 = 8'h1 == _T_21 ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3086 = 8'h2 == _T_21 ? $signed(regsA_2_im) : $signed(_GEN_3085); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3087 = 8'h3 == _T_21 ? $signed(regsA_3_im) : $signed(_GEN_3086); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3088 = 8'h4 == _T_21 ? $signed(regsA_4_im) : $signed(_GEN_3087); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3089 = 8'h5 == _T_21 ? $signed(regsA_5_im) : $signed(_GEN_3088); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3090 = 8'h6 == _T_21 ? $signed(regsA_6_im) : $signed(_GEN_3089); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3091 = 8'h7 == _T_21 ? $signed(regsA_7_im) : $signed(_GEN_3090); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3092 = 8'h8 == _T_21 ? $signed(regsA_8_im) : $signed(_GEN_3091); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3093 = 8'h9 == _T_21 ? $signed(regsA_9_im) : $signed(_GEN_3092); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3094 = 8'ha == _T_21 ? $signed(32'sh0) : $signed(_GEN_3093); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3095 = 8'hb == _T_21 ? $signed(32'sh0) : $signed(_GEN_3094); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3096 = 8'hc == _T_21 ? $signed(32'sh0) : $signed(_GEN_3095); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3097 = 8'hd == _T_21 ? $signed(32'sh0) : $signed(_GEN_3096); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3098 = 8'he == _T_21 ? $signed(32'sh0) : $signed(_GEN_3097); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3099 = 8'hf == _T_21 ? $signed(32'sh0) : $signed(_GEN_3098); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3100 = 8'h10 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3099); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3101 = 8'h11 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3100); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3102 = 8'h12 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3101); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3103 = 8'h13 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3102); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3104 = 8'h14 == _T_21 ? $signed(regsA_10_im) : $signed(_GEN_3103); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3105 = 8'h15 == _T_21 ? $signed(regsA_11_im) : $signed(_GEN_3104); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3106 = 8'h16 == _T_21 ? $signed(regsA_12_im) : $signed(_GEN_3105); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3107 = 8'h17 == _T_21 ? $signed(regsA_13_im) : $signed(_GEN_3106); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3108 = 8'h18 == _T_21 ? $signed(regsA_14_im) : $signed(_GEN_3107); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3109 = 8'h19 == _T_21 ? $signed(regsA_15_im) : $signed(_GEN_3108); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3110 = 8'h1a == _T_21 ? $signed(regsA_16_im) : $signed(_GEN_3109); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3111 = 8'h1b == _T_21 ? $signed(regsA_17_im) : $signed(_GEN_3110); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3112 = 8'h1c == _T_21 ? $signed(regsA_18_im) : $signed(_GEN_3111); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3113 = 8'h1d == _T_21 ? $signed(regsA_19_im) : $signed(_GEN_3112); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3114 = 8'h1e == _T_21 ? $signed(32'sh0) : $signed(_GEN_3113); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3115 = 8'h1f == _T_21 ? $signed(32'sh0) : $signed(_GEN_3114); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3116 = 8'h20 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3115); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3117 = 8'h21 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3116); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3118 = 8'h22 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3117); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3119 = 8'h23 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3118); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3120 = 8'h24 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3119); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3121 = 8'h25 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3120); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3122 = 8'h26 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3121); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3123 = 8'h27 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3122); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3124 = 8'h28 == _T_21 ? $signed(regsA_20_im) : $signed(_GEN_3123); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3125 = 8'h29 == _T_21 ? $signed(regsA_21_im) : $signed(_GEN_3124); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3126 = 8'h2a == _T_21 ? $signed(regsA_22_im) : $signed(_GEN_3125); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3127 = 8'h2b == _T_21 ? $signed(regsA_23_im) : $signed(_GEN_3126); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3128 = 8'h2c == _T_21 ? $signed(regsA_24_im) : $signed(_GEN_3127); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3129 = 8'h2d == _T_21 ? $signed(regsA_25_im) : $signed(_GEN_3128); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3130 = 8'h2e == _T_21 ? $signed(regsA_26_im) : $signed(_GEN_3129); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3131 = 8'h2f == _T_21 ? $signed(regsA_27_im) : $signed(_GEN_3130); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3132 = 8'h30 == _T_21 ? $signed(regsA_28_im) : $signed(_GEN_3131); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3133 = 8'h31 == _T_21 ? $signed(regsA_29_im) : $signed(_GEN_3132); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3134 = 8'h32 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3133); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3135 = 8'h33 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3134); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3136 = 8'h34 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3135); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3137 = 8'h35 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3136); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3138 = 8'h36 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3137); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3139 = 8'h37 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3138); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3140 = 8'h38 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3139); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3141 = 8'h39 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3140); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3142 = 8'h3a == _T_21 ? $signed(32'sh0) : $signed(_GEN_3141); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3143 = 8'h3b == _T_21 ? $signed(32'sh0) : $signed(_GEN_3142); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3144 = 8'h3c == _T_21 ? $signed(regsA_30_im) : $signed(_GEN_3143); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3145 = 8'h3d == _T_21 ? $signed(regsA_31_im) : $signed(_GEN_3144); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3146 = 8'h3e == _T_21 ? $signed(regsA_32_im) : $signed(_GEN_3145); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3147 = 8'h3f == _T_21 ? $signed(regsA_33_im) : $signed(_GEN_3146); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3148 = 8'h40 == _T_21 ? $signed(regsA_34_im) : $signed(_GEN_3147); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3149 = 8'h41 == _T_21 ? $signed(regsA_35_im) : $signed(_GEN_3148); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3150 = 8'h42 == _T_21 ? $signed(regsA_36_im) : $signed(_GEN_3149); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3151 = 8'h43 == _T_21 ? $signed(regsA_37_im) : $signed(_GEN_3150); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3152 = 8'h44 == _T_21 ? $signed(regsA_38_im) : $signed(_GEN_3151); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3153 = 8'h45 == _T_21 ? $signed(regsA_39_im) : $signed(_GEN_3152); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3154 = 8'h46 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3153); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3155 = 8'h47 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3154); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3156 = 8'h48 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3155); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3157 = 8'h49 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3156); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3158 = 8'h4a == _T_21 ? $signed(32'sh0) : $signed(_GEN_3157); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3159 = 8'h4b == _T_21 ? $signed(32'sh0) : $signed(_GEN_3158); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3160 = 8'h4c == _T_21 ? $signed(32'sh0) : $signed(_GEN_3159); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3161 = 8'h4d == _T_21 ? $signed(32'sh0) : $signed(_GEN_3160); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3162 = 8'h4e == _T_21 ? $signed(32'sh0) : $signed(_GEN_3161); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3163 = 8'h4f == _T_21 ? $signed(32'sh0) : $signed(_GEN_3162); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3164 = 8'h50 == _T_21 ? $signed(regsA_40_im) : $signed(_GEN_3163); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3165 = 8'h51 == _T_21 ? $signed(regsA_41_im) : $signed(_GEN_3164); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3166 = 8'h52 == _T_21 ? $signed(regsA_42_im) : $signed(_GEN_3165); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3167 = 8'h53 == _T_21 ? $signed(regsA_43_im) : $signed(_GEN_3166); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3168 = 8'h54 == _T_21 ? $signed(regsA_44_im) : $signed(_GEN_3167); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3169 = 8'h55 == _T_21 ? $signed(regsA_45_im) : $signed(_GEN_3168); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3170 = 8'h56 == _T_21 ? $signed(regsA_46_im) : $signed(_GEN_3169); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3171 = 8'h57 == _T_21 ? $signed(regsA_47_im) : $signed(_GEN_3170); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3172 = 8'h58 == _T_21 ? $signed(regsA_48_im) : $signed(_GEN_3171); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3173 = 8'h59 == _T_21 ? $signed(regsA_49_im) : $signed(_GEN_3172); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3174 = 8'h5a == _T_21 ? $signed(32'sh0) : $signed(_GEN_3173); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3175 = 8'h5b == _T_21 ? $signed(32'sh0) : $signed(_GEN_3174); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3176 = 8'h5c == _T_21 ? $signed(32'sh0) : $signed(_GEN_3175); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3177 = 8'h5d == _T_21 ? $signed(32'sh0) : $signed(_GEN_3176); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3178 = 8'h5e == _T_21 ? $signed(32'sh0) : $signed(_GEN_3177); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3179 = 8'h5f == _T_21 ? $signed(32'sh0) : $signed(_GEN_3178); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3180 = 8'h60 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3179); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3181 = 8'h61 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3180); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3182 = 8'h62 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3181); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3183 = 8'h63 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3182); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3184 = 8'h64 == _T_21 ? $signed(regsA_50_im) : $signed(_GEN_3183); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3185 = 8'h65 == _T_21 ? $signed(regsA_51_im) : $signed(_GEN_3184); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3186 = 8'h66 == _T_21 ? $signed(regsA_52_im) : $signed(_GEN_3185); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3187 = 8'h67 == _T_21 ? $signed(regsA_53_im) : $signed(_GEN_3186); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3188 = 8'h68 == _T_21 ? $signed(regsA_54_im) : $signed(_GEN_3187); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3189 = 8'h69 == _T_21 ? $signed(regsA_55_im) : $signed(_GEN_3188); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3190 = 8'h6a == _T_21 ? $signed(regsA_56_im) : $signed(_GEN_3189); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3191 = 8'h6b == _T_21 ? $signed(regsA_57_im) : $signed(_GEN_3190); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3192 = 8'h6c == _T_21 ? $signed(regsA_58_im) : $signed(_GEN_3191); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3193 = 8'h6d == _T_21 ? $signed(regsA_59_im) : $signed(_GEN_3192); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3194 = 8'h6e == _T_21 ? $signed(32'sh0) : $signed(_GEN_3193); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3195 = 8'h6f == _T_21 ? $signed(32'sh0) : $signed(_GEN_3194); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3196 = 8'h70 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3195); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3197 = 8'h71 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3196); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3198 = 8'h72 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3197); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3199 = 8'h73 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3198); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3200 = 8'h74 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3199); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3201 = 8'h75 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3200); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3202 = 8'h76 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3201); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3203 = 8'h77 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3202); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3204 = 8'h78 == _T_21 ? $signed(regsA_60_im) : $signed(_GEN_3203); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3205 = 8'h79 == _T_21 ? $signed(regsA_61_im) : $signed(_GEN_3204); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3206 = 8'h7a == _T_21 ? $signed(regsA_62_im) : $signed(_GEN_3205); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3207 = 8'h7b == _T_21 ? $signed(regsA_63_im) : $signed(_GEN_3206); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3208 = 8'h7c == _T_21 ? $signed(regsA_64_im) : $signed(_GEN_3207); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3209 = 8'h7d == _T_21 ? $signed(regsA_65_im) : $signed(_GEN_3208); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3210 = 8'h7e == _T_21 ? $signed(regsA_66_im) : $signed(_GEN_3209); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3211 = 8'h7f == _T_21 ? $signed(regsA_67_im) : $signed(_GEN_3210); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3212 = 8'h80 == _T_21 ? $signed(regsA_68_im) : $signed(_GEN_3211); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3213 = 8'h81 == _T_21 ? $signed(regsA_69_im) : $signed(_GEN_3212); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3214 = 8'h82 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3213); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3215 = 8'h83 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3214); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3216 = 8'h84 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3215); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3217 = 8'h85 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3216); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3218 = 8'h86 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3217); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3219 = 8'h87 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3218); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3220 = 8'h88 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3219); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3221 = 8'h89 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3220); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3222 = 8'h8a == _T_21 ? $signed(32'sh0) : $signed(_GEN_3221); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3223 = 8'h8b == _T_21 ? $signed(32'sh0) : $signed(_GEN_3222); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3224 = 8'h8c == _T_21 ? $signed(regsA_70_im) : $signed(_GEN_3223); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3225 = 8'h8d == _T_21 ? $signed(regsA_71_im) : $signed(_GEN_3224); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3226 = 8'h8e == _T_21 ? $signed(regsA_72_im) : $signed(_GEN_3225); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3227 = 8'h8f == _T_21 ? $signed(regsA_73_im) : $signed(_GEN_3226); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3228 = 8'h90 == _T_21 ? $signed(regsA_74_im) : $signed(_GEN_3227); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3229 = 8'h91 == _T_21 ? $signed(regsA_75_im) : $signed(_GEN_3228); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3230 = 8'h92 == _T_21 ? $signed(regsA_76_im) : $signed(_GEN_3229); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3231 = 8'h93 == _T_21 ? $signed(regsA_77_im) : $signed(_GEN_3230); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3232 = 8'h94 == _T_21 ? $signed(regsA_78_im) : $signed(_GEN_3231); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3233 = 8'h95 == _T_21 ? $signed(regsA_79_im) : $signed(_GEN_3232); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3234 = 8'h96 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3233); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3235 = 8'h97 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3234); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3236 = 8'h98 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3235); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3237 = 8'h99 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3236); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3238 = 8'h9a == _T_21 ? $signed(32'sh0) : $signed(_GEN_3237); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3239 = 8'h9b == _T_21 ? $signed(32'sh0) : $signed(_GEN_3238); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3240 = 8'h9c == _T_21 ? $signed(32'sh0) : $signed(_GEN_3239); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3241 = 8'h9d == _T_21 ? $signed(32'sh0) : $signed(_GEN_3240); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3242 = 8'h9e == _T_21 ? $signed(32'sh0) : $signed(_GEN_3241); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3243 = 8'h9f == _T_21 ? $signed(32'sh0) : $signed(_GEN_3242); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3244 = 8'ha0 == _T_21 ? $signed(regsA_80_im) : $signed(_GEN_3243); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3245 = 8'ha1 == _T_21 ? $signed(regsA_81_im) : $signed(_GEN_3244); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3246 = 8'ha2 == _T_21 ? $signed(regsA_82_im) : $signed(_GEN_3245); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3247 = 8'ha3 == _T_21 ? $signed(regsA_83_im) : $signed(_GEN_3246); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3248 = 8'ha4 == _T_21 ? $signed(regsA_84_im) : $signed(_GEN_3247); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3249 = 8'ha5 == _T_21 ? $signed(regsA_85_im) : $signed(_GEN_3248); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3250 = 8'ha6 == _T_21 ? $signed(regsA_86_im) : $signed(_GEN_3249); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3251 = 8'ha7 == _T_21 ? $signed(regsA_87_im) : $signed(_GEN_3250); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3252 = 8'ha8 == _T_21 ? $signed(regsA_88_im) : $signed(_GEN_3251); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3253 = 8'ha9 == _T_21 ? $signed(regsA_89_im) : $signed(_GEN_3252); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3254 = 8'haa == _T_21 ? $signed(32'sh0) : $signed(_GEN_3253); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3255 = 8'hab == _T_21 ? $signed(32'sh0) : $signed(_GEN_3254); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3256 = 8'hac == _T_21 ? $signed(32'sh0) : $signed(_GEN_3255); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3257 = 8'had == _T_21 ? $signed(32'sh0) : $signed(_GEN_3256); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3258 = 8'hae == _T_21 ? $signed(32'sh0) : $signed(_GEN_3257); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3259 = 8'haf == _T_21 ? $signed(32'sh0) : $signed(_GEN_3258); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3260 = 8'hb0 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3259); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3261 = 8'hb1 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3260); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3262 = 8'hb2 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3261); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3263 = 8'hb3 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3262); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3264 = 8'hb4 == _T_21 ? $signed(regsA_90_im) : $signed(_GEN_3263); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3265 = 8'hb5 == _T_21 ? $signed(regsA_91_im) : $signed(_GEN_3264); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3266 = 8'hb6 == _T_21 ? $signed(regsA_92_im) : $signed(_GEN_3265); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3267 = 8'hb7 == _T_21 ? $signed(regsA_93_im) : $signed(_GEN_3266); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3268 = 8'hb8 == _T_21 ? $signed(regsA_94_im) : $signed(_GEN_3267); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3269 = 8'hb9 == _T_21 ? $signed(regsA_95_im) : $signed(_GEN_3268); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3270 = 8'hba == _T_21 ? $signed(regsA_96_im) : $signed(_GEN_3269); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3271 = 8'hbb == _T_21 ? $signed(regsA_97_im) : $signed(_GEN_3270); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3272 = 8'hbc == _T_21 ? $signed(regsA_98_im) : $signed(_GEN_3271); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3273 = 8'hbd == _T_21 ? $signed(regsA_99_im) : $signed(_GEN_3272); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3275 = 8'h1 == _T_21 ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3276 = 8'h2 == _T_21 ? $signed(regsA_2_re) : $signed(_GEN_3275); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3277 = 8'h3 == _T_21 ? $signed(regsA_3_re) : $signed(_GEN_3276); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3278 = 8'h4 == _T_21 ? $signed(regsA_4_re) : $signed(_GEN_3277); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3279 = 8'h5 == _T_21 ? $signed(regsA_5_re) : $signed(_GEN_3278); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3280 = 8'h6 == _T_21 ? $signed(regsA_6_re) : $signed(_GEN_3279); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3281 = 8'h7 == _T_21 ? $signed(regsA_7_re) : $signed(_GEN_3280); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3282 = 8'h8 == _T_21 ? $signed(regsA_8_re) : $signed(_GEN_3281); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3283 = 8'h9 == _T_21 ? $signed(regsA_9_re) : $signed(_GEN_3282); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3284 = 8'ha == _T_21 ? $signed(32'sh0) : $signed(_GEN_3283); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3285 = 8'hb == _T_21 ? $signed(32'sh0) : $signed(_GEN_3284); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3286 = 8'hc == _T_21 ? $signed(32'sh0) : $signed(_GEN_3285); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3287 = 8'hd == _T_21 ? $signed(32'sh0) : $signed(_GEN_3286); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3288 = 8'he == _T_21 ? $signed(32'sh0) : $signed(_GEN_3287); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3289 = 8'hf == _T_21 ? $signed(32'sh0) : $signed(_GEN_3288); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3290 = 8'h10 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3289); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3291 = 8'h11 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3290); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3292 = 8'h12 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3291); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3293 = 8'h13 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3292); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3294 = 8'h14 == _T_21 ? $signed(regsA_10_re) : $signed(_GEN_3293); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3295 = 8'h15 == _T_21 ? $signed(regsA_11_re) : $signed(_GEN_3294); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3296 = 8'h16 == _T_21 ? $signed(regsA_12_re) : $signed(_GEN_3295); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3297 = 8'h17 == _T_21 ? $signed(regsA_13_re) : $signed(_GEN_3296); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3298 = 8'h18 == _T_21 ? $signed(regsA_14_re) : $signed(_GEN_3297); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3299 = 8'h19 == _T_21 ? $signed(regsA_15_re) : $signed(_GEN_3298); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3300 = 8'h1a == _T_21 ? $signed(regsA_16_re) : $signed(_GEN_3299); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3301 = 8'h1b == _T_21 ? $signed(regsA_17_re) : $signed(_GEN_3300); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3302 = 8'h1c == _T_21 ? $signed(regsA_18_re) : $signed(_GEN_3301); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3303 = 8'h1d == _T_21 ? $signed(regsA_19_re) : $signed(_GEN_3302); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3304 = 8'h1e == _T_21 ? $signed(32'sh0) : $signed(_GEN_3303); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3305 = 8'h1f == _T_21 ? $signed(32'sh0) : $signed(_GEN_3304); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3306 = 8'h20 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3305); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3307 = 8'h21 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3306); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3308 = 8'h22 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3307); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3309 = 8'h23 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3308); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3310 = 8'h24 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3309); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3311 = 8'h25 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3310); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3312 = 8'h26 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3311); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3313 = 8'h27 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3312); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3314 = 8'h28 == _T_21 ? $signed(regsA_20_re) : $signed(_GEN_3313); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3315 = 8'h29 == _T_21 ? $signed(regsA_21_re) : $signed(_GEN_3314); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3316 = 8'h2a == _T_21 ? $signed(regsA_22_re) : $signed(_GEN_3315); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3317 = 8'h2b == _T_21 ? $signed(regsA_23_re) : $signed(_GEN_3316); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3318 = 8'h2c == _T_21 ? $signed(regsA_24_re) : $signed(_GEN_3317); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3319 = 8'h2d == _T_21 ? $signed(regsA_25_re) : $signed(_GEN_3318); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3320 = 8'h2e == _T_21 ? $signed(regsA_26_re) : $signed(_GEN_3319); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3321 = 8'h2f == _T_21 ? $signed(regsA_27_re) : $signed(_GEN_3320); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3322 = 8'h30 == _T_21 ? $signed(regsA_28_re) : $signed(_GEN_3321); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3323 = 8'h31 == _T_21 ? $signed(regsA_29_re) : $signed(_GEN_3322); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3324 = 8'h32 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3323); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3325 = 8'h33 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3324); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3326 = 8'h34 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3325); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3327 = 8'h35 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3326); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3328 = 8'h36 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3327); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3329 = 8'h37 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3328); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3330 = 8'h38 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3329); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3331 = 8'h39 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3330); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3332 = 8'h3a == _T_21 ? $signed(32'sh0) : $signed(_GEN_3331); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3333 = 8'h3b == _T_21 ? $signed(32'sh0) : $signed(_GEN_3332); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3334 = 8'h3c == _T_21 ? $signed(regsA_30_re) : $signed(_GEN_3333); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3335 = 8'h3d == _T_21 ? $signed(regsA_31_re) : $signed(_GEN_3334); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3336 = 8'h3e == _T_21 ? $signed(regsA_32_re) : $signed(_GEN_3335); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3337 = 8'h3f == _T_21 ? $signed(regsA_33_re) : $signed(_GEN_3336); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3338 = 8'h40 == _T_21 ? $signed(regsA_34_re) : $signed(_GEN_3337); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3339 = 8'h41 == _T_21 ? $signed(regsA_35_re) : $signed(_GEN_3338); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3340 = 8'h42 == _T_21 ? $signed(regsA_36_re) : $signed(_GEN_3339); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3341 = 8'h43 == _T_21 ? $signed(regsA_37_re) : $signed(_GEN_3340); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3342 = 8'h44 == _T_21 ? $signed(regsA_38_re) : $signed(_GEN_3341); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3343 = 8'h45 == _T_21 ? $signed(regsA_39_re) : $signed(_GEN_3342); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3344 = 8'h46 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3343); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3345 = 8'h47 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3344); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3346 = 8'h48 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3345); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3347 = 8'h49 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3346); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3348 = 8'h4a == _T_21 ? $signed(32'sh0) : $signed(_GEN_3347); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3349 = 8'h4b == _T_21 ? $signed(32'sh0) : $signed(_GEN_3348); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3350 = 8'h4c == _T_21 ? $signed(32'sh0) : $signed(_GEN_3349); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3351 = 8'h4d == _T_21 ? $signed(32'sh0) : $signed(_GEN_3350); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3352 = 8'h4e == _T_21 ? $signed(32'sh0) : $signed(_GEN_3351); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3353 = 8'h4f == _T_21 ? $signed(32'sh0) : $signed(_GEN_3352); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3354 = 8'h50 == _T_21 ? $signed(regsA_40_re) : $signed(_GEN_3353); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3355 = 8'h51 == _T_21 ? $signed(regsA_41_re) : $signed(_GEN_3354); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3356 = 8'h52 == _T_21 ? $signed(regsA_42_re) : $signed(_GEN_3355); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3357 = 8'h53 == _T_21 ? $signed(regsA_43_re) : $signed(_GEN_3356); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3358 = 8'h54 == _T_21 ? $signed(regsA_44_re) : $signed(_GEN_3357); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3359 = 8'h55 == _T_21 ? $signed(regsA_45_re) : $signed(_GEN_3358); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3360 = 8'h56 == _T_21 ? $signed(regsA_46_re) : $signed(_GEN_3359); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3361 = 8'h57 == _T_21 ? $signed(regsA_47_re) : $signed(_GEN_3360); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3362 = 8'h58 == _T_21 ? $signed(regsA_48_re) : $signed(_GEN_3361); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3363 = 8'h59 == _T_21 ? $signed(regsA_49_re) : $signed(_GEN_3362); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3364 = 8'h5a == _T_21 ? $signed(32'sh0) : $signed(_GEN_3363); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3365 = 8'h5b == _T_21 ? $signed(32'sh0) : $signed(_GEN_3364); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3366 = 8'h5c == _T_21 ? $signed(32'sh0) : $signed(_GEN_3365); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3367 = 8'h5d == _T_21 ? $signed(32'sh0) : $signed(_GEN_3366); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3368 = 8'h5e == _T_21 ? $signed(32'sh0) : $signed(_GEN_3367); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3369 = 8'h5f == _T_21 ? $signed(32'sh0) : $signed(_GEN_3368); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3370 = 8'h60 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3369); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3371 = 8'h61 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3370); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3372 = 8'h62 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3371); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3373 = 8'h63 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3372); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3374 = 8'h64 == _T_21 ? $signed(regsA_50_re) : $signed(_GEN_3373); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3375 = 8'h65 == _T_21 ? $signed(regsA_51_re) : $signed(_GEN_3374); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3376 = 8'h66 == _T_21 ? $signed(regsA_52_re) : $signed(_GEN_3375); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3377 = 8'h67 == _T_21 ? $signed(regsA_53_re) : $signed(_GEN_3376); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3378 = 8'h68 == _T_21 ? $signed(regsA_54_re) : $signed(_GEN_3377); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3379 = 8'h69 == _T_21 ? $signed(regsA_55_re) : $signed(_GEN_3378); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3380 = 8'h6a == _T_21 ? $signed(regsA_56_re) : $signed(_GEN_3379); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3381 = 8'h6b == _T_21 ? $signed(regsA_57_re) : $signed(_GEN_3380); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3382 = 8'h6c == _T_21 ? $signed(regsA_58_re) : $signed(_GEN_3381); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3383 = 8'h6d == _T_21 ? $signed(regsA_59_re) : $signed(_GEN_3382); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3384 = 8'h6e == _T_21 ? $signed(32'sh0) : $signed(_GEN_3383); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3385 = 8'h6f == _T_21 ? $signed(32'sh0) : $signed(_GEN_3384); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3386 = 8'h70 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3385); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3387 = 8'h71 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3386); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3388 = 8'h72 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3387); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3389 = 8'h73 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3388); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3390 = 8'h74 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3389); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3391 = 8'h75 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3390); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3392 = 8'h76 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3391); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3393 = 8'h77 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3392); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3394 = 8'h78 == _T_21 ? $signed(regsA_60_re) : $signed(_GEN_3393); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3395 = 8'h79 == _T_21 ? $signed(regsA_61_re) : $signed(_GEN_3394); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3396 = 8'h7a == _T_21 ? $signed(regsA_62_re) : $signed(_GEN_3395); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3397 = 8'h7b == _T_21 ? $signed(regsA_63_re) : $signed(_GEN_3396); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3398 = 8'h7c == _T_21 ? $signed(regsA_64_re) : $signed(_GEN_3397); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3399 = 8'h7d == _T_21 ? $signed(regsA_65_re) : $signed(_GEN_3398); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3400 = 8'h7e == _T_21 ? $signed(regsA_66_re) : $signed(_GEN_3399); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3401 = 8'h7f == _T_21 ? $signed(regsA_67_re) : $signed(_GEN_3400); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3402 = 8'h80 == _T_21 ? $signed(regsA_68_re) : $signed(_GEN_3401); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3403 = 8'h81 == _T_21 ? $signed(regsA_69_re) : $signed(_GEN_3402); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3404 = 8'h82 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3403); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3405 = 8'h83 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3404); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3406 = 8'h84 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3405); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3407 = 8'h85 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3406); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3408 = 8'h86 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3407); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3409 = 8'h87 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3408); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3410 = 8'h88 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3409); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3411 = 8'h89 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3410); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3412 = 8'h8a == _T_21 ? $signed(32'sh0) : $signed(_GEN_3411); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3413 = 8'h8b == _T_21 ? $signed(32'sh0) : $signed(_GEN_3412); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3414 = 8'h8c == _T_21 ? $signed(regsA_70_re) : $signed(_GEN_3413); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3415 = 8'h8d == _T_21 ? $signed(regsA_71_re) : $signed(_GEN_3414); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3416 = 8'h8e == _T_21 ? $signed(regsA_72_re) : $signed(_GEN_3415); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3417 = 8'h8f == _T_21 ? $signed(regsA_73_re) : $signed(_GEN_3416); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3418 = 8'h90 == _T_21 ? $signed(regsA_74_re) : $signed(_GEN_3417); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3419 = 8'h91 == _T_21 ? $signed(regsA_75_re) : $signed(_GEN_3418); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3420 = 8'h92 == _T_21 ? $signed(regsA_76_re) : $signed(_GEN_3419); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3421 = 8'h93 == _T_21 ? $signed(regsA_77_re) : $signed(_GEN_3420); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3422 = 8'h94 == _T_21 ? $signed(regsA_78_re) : $signed(_GEN_3421); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3423 = 8'h95 == _T_21 ? $signed(regsA_79_re) : $signed(_GEN_3422); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3424 = 8'h96 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3423); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3425 = 8'h97 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3424); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3426 = 8'h98 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3425); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3427 = 8'h99 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3426); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3428 = 8'h9a == _T_21 ? $signed(32'sh0) : $signed(_GEN_3427); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3429 = 8'h9b == _T_21 ? $signed(32'sh0) : $signed(_GEN_3428); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3430 = 8'h9c == _T_21 ? $signed(32'sh0) : $signed(_GEN_3429); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3431 = 8'h9d == _T_21 ? $signed(32'sh0) : $signed(_GEN_3430); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3432 = 8'h9e == _T_21 ? $signed(32'sh0) : $signed(_GEN_3431); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3433 = 8'h9f == _T_21 ? $signed(32'sh0) : $signed(_GEN_3432); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3434 = 8'ha0 == _T_21 ? $signed(regsA_80_re) : $signed(_GEN_3433); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3435 = 8'ha1 == _T_21 ? $signed(regsA_81_re) : $signed(_GEN_3434); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3436 = 8'ha2 == _T_21 ? $signed(regsA_82_re) : $signed(_GEN_3435); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3437 = 8'ha3 == _T_21 ? $signed(regsA_83_re) : $signed(_GEN_3436); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3438 = 8'ha4 == _T_21 ? $signed(regsA_84_re) : $signed(_GEN_3437); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3439 = 8'ha5 == _T_21 ? $signed(regsA_85_re) : $signed(_GEN_3438); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3440 = 8'ha6 == _T_21 ? $signed(regsA_86_re) : $signed(_GEN_3439); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3441 = 8'ha7 == _T_21 ? $signed(regsA_87_re) : $signed(_GEN_3440); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3442 = 8'ha8 == _T_21 ? $signed(regsA_88_re) : $signed(_GEN_3441); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3443 = 8'ha9 == _T_21 ? $signed(regsA_89_re) : $signed(_GEN_3442); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3444 = 8'haa == _T_21 ? $signed(32'sh0) : $signed(_GEN_3443); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3445 = 8'hab == _T_21 ? $signed(32'sh0) : $signed(_GEN_3444); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3446 = 8'hac == _T_21 ? $signed(32'sh0) : $signed(_GEN_3445); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3447 = 8'had == _T_21 ? $signed(32'sh0) : $signed(_GEN_3446); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3448 = 8'hae == _T_21 ? $signed(32'sh0) : $signed(_GEN_3447); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3449 = 8'haf == _T_21 ? $signed(32'sh0) : $signed(_GEN_3448); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3450 = 8'hb0 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3449); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3451 = 8'hb1 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3450); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3452 = 8'hb2 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3451); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3453 = 8'hb3 == _T_21 ? $signed(32'sh0) : $signed(_GEN_3452); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3454 = 8'hb4 == _T_21 ? $signed(regsA_90_re) : $signed(_GEN_3453); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3455 = 8'hb5 == _T_21 ? $signed(regsA_91_re) : $signed(_GEN_3454); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3456 = 8'hb6 == _T_21 ? $signed(regsA_92_re) : $signed(_GEN_3455); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3457 = 8'hb7 == _T_21 ? $signed(regsA_93_re) : $signed(_GEN_3456); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3458 = 8'hb8 == _T_21 ? $signed(regsA_94_re) : $signed(_GEN_3457); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3459 = 8'hb9 == _T_21 ? $signed(regsA_95_re) : $signed(_GEN_3458); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3460 = 8'hba == _T_21 ? $signed(regsA_96_re) : $signed(_GEN_3459); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3461 = 8'hbb == _T_21 ? $signed(regsA_97_re) : $signed(_GEN_3460); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3462 = 8'hbc == _T_21 ? $signed(regsA_98_re) : $signed(_GEN_3461); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3463 = 8'hbd == _T_21 ? $signed(regsA_99_re) : $signed(_GEN_3462); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [7:0] _T_22 = 3'h7 * 5'h13; // @[Matrix_Mul_V1.scala 148:44]
  wire [7:0] _T_24 = _T_22 + _GEN_9199; // @[Matrix_Mul_V1.scala 148:60]
  wire [31:0] _GEN_3465 = 8'h1 == _T_24 ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3466 = 8'h2 == _T_24 ? $signed(regsA_2_im) : $signed(_GEN_3465); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3467 = 8'h3 == _T_24 ? $signed(regsA_3_im) : $signed(_GEN_3466); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3468 = 8'h4 == _T_24 ? $signed(regsA_4_im) : $signed(_GEN_3467); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3469 = 8'h5 == _T_24 ? $signed(regsA_5_im) : $signed(_GEN_3468); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3470 = 8'h6 == _T_24 ? $signed(regsA_6_im) : $signed(_GEN_3469); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3471 = 8'h7 == _T_24 ? $signed(regsA_7_im) : $signed(_GEN_3470); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3472 = 8'h8 == _T_24 ? $signed(regsA_8_im) : $signed(_GEN_3471); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3473 = 8'h9 == _T_24 ? $signed(regsA_9_im) : $signed(_GEN_3472); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3474 = 8'ha == _T_24 ? $signed(32'sh0) : $signed(_GEN_3473); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3475 = 8'hb == _T_24 ? $signed(32'sh0) : $signed(_GEN_3474); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3476 = 8'hc == _T_24 ? $signed(32'sh0) : $signed(_GEN_3475); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3477 = 8'hd == _T_24 ? $signed(32'sh0) : $signed(_GEN_3476); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3478 = 8'he == _T_24 ? $signed(32'sh0) : $signed(_GEN_3477); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3479 = 8'hf == _T_24 ? $signed(32'sh0) : $signed(_GEN_3478); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3480 = 8'h10 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3479); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3481 = 8'h11 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3480); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3482 = 8'h12 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3481); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3483 = 8'h13 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3482); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3484 = 8'h14 == _T_24 ? $signed(regsA_10_im) : $signed(_GEN_3483); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3485 = 8'h15 == _T_24 ? $signed(regsA_11_im) : $signed(_GEN_3484); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3486 = 8'h16 == _T_24 ? $signed(regsA_12_im) : $signed(_GEN_3485); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3487 = 8'h17 == _T_24 ? $signed(regsA_13_im) : $signed(_GEN_3486); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3488 = 8'h18 == _T_24 ? $signed(regsA_14_im) : $signed(_GEN_3487); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3489 = 8'h19 == _T_24 ? $signed(regsA_15_im) : $signed(_GEN_3488); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3490 = 8'h1a == _T_24 ? $signed(regsA_16_im) : $signed(_GEN_3489); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3491 = 8'h1b == _T_24 ? $signed(regsA_17_im) : $signed(_GEN_3490); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3492 = 8'h1c == _T_24 ? $signed(regsA_18_im) : $signed(_GEN_3491); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3493 = 8'h1d == _T_24 ? $signed(regsA_19_im) : $signed(_GEN_3492); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3494 = 8'h1e == _T_24 ? $signed(32'sh0) : $signed(_GEN_3493); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3495 = 8'h1f == _T_24 ? $signed(32'sh0) : $signed(_GEN_3494); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3496 = 8'h20 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3495); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3497 = 8'h21 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3496); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3498 = 8'h22 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3497); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3499 = 8'h23 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3498); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3500 = 8'h24 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3499); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3501 = 8'h25 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3500); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3502 = 8'h26 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3501); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3503 = 8'h27 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3502); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3504 = 8'h28 == _T_24 ? $signed(regsA_20_im) : $signed(_GEN_3503); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3505 = 8'h29 == _T_24 ? $signed(regsA_21_im) : $signed(_GEN_3504); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3506 = 8'h2a == _T_24 ? $signed(regsA_22_im) : $signed(_GEN_3505); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3507 = 8'h2b == _T_24 ? $signed(regsA_23_im) : $signed(_GEN_3506); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3508 = 8'h2c == _T_24 ? $signed(regsA_24_im) : $signed(_GEN_3507); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3509 = 8'h2d == _T_24 ? $signed(regsA_25_im) : $signed(_GEN_3508); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3510 = 8'h2e == _T_24 ? $signed(regsA_26_im) : $signed(_GEN_3509); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3511 = 8'h2f == _T_24 ? $signed(regsA_27_im) : $signed(_GEN_3510); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3512 = 8'h30 == _T_24 ? $signed(regsA_28_im) : $signed(_GEN_3511); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3513 = 8'h31 == _T_24 ? $signed(regsA_29_im) : $signed(_GEN_3512); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3514 = 8'h32 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3513); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3515 = 8'h33 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3514); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3516 = 8'h34 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3515); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3517 = 8'h35 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3516); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3518 = 8'h36 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3517); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3519 = 8'h37 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3518); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3520 = 8'h38 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3519); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3521 = 8'h39 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3520); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3522 = 8'h3a == _T_24 ? $signed(32'sh0) : $signed(_GEN_3521); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3523 = 8'h3b == _T_24 ? $signed(32'sh0) : $signed(_GEN_3522); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3524 = 8'h3c == _T_24 ? $signed(regsA_30_im) : $signed(_GEN_3523); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3525 = 8'h3d == _T_24 ? $signed(regsA_31_im) : $signed(_GEN_3524); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3526 = 8'h3e == _T_24 ? $signed(regsA_32_im) : $signed(_GEN_3525); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3527 = 8'h3f == _T_24 ? $signed(regsA_33_im) : $signed(_GEN_3526); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3528 = 8'h40 == _T_24 ? $signed(regsA_34_im) : $signed(_GEN_3527); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3529 = 8'h41 == _T_24 ? $signed(regsA_35_im) : $signed(_GEN_3528); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3530 = 8'h42 == _T_24 ? $signed(regsA_36_im) : $signed(_GEN_3529); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3531 = 8'h43 == _T_24 ? $signed(regsA_37_im) : $signed(_GEN_3530); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3532 = 8'h44 == _T_24 ? $signed(regsA_38_im) : $signed(_GEN_3531); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3533 = 8'h45 == _T_24 ? $signed(regsA_39_im) : $signed(_GEN_3532); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3534 = 8'h46 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3533); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3535 = 8'h47 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3534); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3536 = 8'h48 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3535); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3537 = 8'h49 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3536); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3538 = 8'h4a == _T_24 ? $signed(32'sh0) : $signed(_GEN_3537); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3539 = 8'h4b == _T_24 ? $signed(32'sh0) : $signed(_GEN_3538); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3540 = 8'h4c == _T_24 ? $signed(32'sh0) : $signed(_GEN_3539); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3541 = 8'h4d == _T_24 ? $signed(32'sh0) : $signed(_GEN_3540); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3542 = 8'h4e == _T_24 ? $signed(32'sh0) : $signed(_GEN_3541); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3543 = 8'h4f == _T_24 ? $signed(32'sh0) : $signed(_GEN_3542); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3544 = 8'h50 == _T_24 ? $signed(regsA_40_im) : $signed(_GEN_3543); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3545 = 8'h51 == _T_24 ? $signed(regsA_41_im) : $signed(_GEN_3544); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3546 = 8'h52 == _T_24 ? $signed(regsA_42_im) : $signed(_GEN_3545); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3547 = 8'h53 == _T_24 ? $signed(regsA_43_im) : $signed(_GEN_3546); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3548 = 8'h54 == _T_24 ? $signed(regsA_44_im) : $signed(_GEN_3547); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3549 = 8'h55 == _T_24 ? $signed(regsA_45_im) : $signed(_GEN_3548); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3550 = 8'h56 == _T_24 ? $signed(regsA_46_im) : $signed(_GEN_3549); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3551 = 8'h57 == _T_24 ? $signed(regsA_47_im) : $signed(_GEN_3550); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3552 = 8'h58 == _T_24 ? $signed(regsA_48_im) : $signed(_GEN_3551); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3553 = 8'h59 == _T_24 ? $signed(regsA_49_im) : $signed(_GEN_3552); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3554 = 8'h5a == _T_24 ? $signed(32'sh0) : $signed(_GEN_3553); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3555 = 8'h5b == _T_24 ? $signed(32'sh0) : $signed(_GEN_3554); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3556 = 8'h5c == _T_24 ? $signed(32'sh0) : $signed(_GEN_3555); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3557 = 8'h5d == _T_24 ? $signed(32'sh0) : $signed(_GEN_3556); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3558 = 8'h5e == _T_24 ? $signed(32'sh0) : $signed(_GEN_3557); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3559 = 8'h5f == _T_24 ? $signed(32'sh0) : $signed(_GEN_3558); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3560 = 8'h60 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3559); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3561 = 8'h61 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3560); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3562 = 8'h62 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3561); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3563 = 8'h63 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3562); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3564 = 8'h64 == _T_24 ? $signed(regsA_50_im) : $signed(_GEN_3563); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3565 = 8'h65 == _T_24 ? $signed(regsA_51_im) : $signed(_GEN_3564); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3566 = 8'h66 == _T_24 ? $signed(regsA_52_im) : $signed(_GEN_3565); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3567 = 8'h67 == _T_24 ? $signed(regsA_53_im) : $signed(_GEN_3566); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3568 = 8'h68 == _T_24 ? $signed(regsA_54_im) : $signed(_GEN_3567); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3569 = 8'h69 == _T_24 ? $signed(regsA_55_im) : $signed(_GEN_3568); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3570 = 8'h6a == _T_24 ? $signed(regsA_56_im) : $signed(_GEN_3569); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3571 = 8'h6b == _T_24 ? $signed(regsA_57_im) : $signed(_GEN_3570); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3572 = 8'h6c == _T_24 ? $signed(regsA_58_im) : $signed(_GEN_3571); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3573 = 8'h6d == _T_24 ? $signed(regsA_59_im) : $signed(_GEN_3572); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3574 = 8'h6e == _T_24 ? $signed(32'sh0) : $signed(_GEN_3573); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3575 = 8'h6f == _T_24 ? $signed(32'sh0) : $signed(_GEN_3574); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3576 = 8'h70 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3575); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3577 = 8'h71 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3576); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3578 = 8'h72 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3577); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3579 = 8'h73 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3578); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3580 = 8'h74 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3579); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3581 = 8'h75 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3580); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3582 = 8'h76 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3581); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3583 = 8'h77 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3582); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3584 = 8'h78 == _T_24 ? $signed(regsA_60_im) : $signed(_GEN_3583); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3585 = 8'h79 == _T_24 ? $signed(regsA_61_im) : $signed(_GEN_3584); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3586 = 8'h7a == _T_24 ? $signed(regsA_62_im) : $signed(_GEN_3585); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3587 = 8'h7b == _T_24 ? $signed(regsA_63_im) : $signed(_GEN_3586); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3588 = 8'h7c == _T_24 ? $signed(regsA_64_im) : $signed(_GEN_3587); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3589 = 8'h7d == _T_24 ? $signed(regsA_65_im) : $signed(_GEN_3588); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3590 = 8'h7e == _T_24 ? $signed(regsA_66_im) : $signed(_GEN_3589); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3591 = 8'h7f == _T_24 ? $signed(regsA_67_im) : $signed(_GEN_3590); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3592 = 8'h80 == _T_24 ? $signed(regsA_68_im) : $signed(_GEN_3591); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3593 = 8'h81 == _T_24 ? $signed(regsA_69_im) : $signed(_GEN_3592); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3594 = 8'h82 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3593); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3595 = 8'h83 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3594); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3596 = 8'h84 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3595); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3597 = 8'h85 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3596); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3598 = 8'h86 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3597); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3599 = 8'h87 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3598); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3600 = 8'h88 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3599); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3601 = 8'h89 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3600); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3602 = 8'h8a == _T_24 ? $signed(32'sh0) : $signed(_GEN_3601); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3603 = 8'h8b == _T_24 ? $signed(32'sh0) : $signed(_GEN_3602); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3604 = 8'h8c == _T_24 ? $signed(regsA_70_im) : $signed(_GEN_3603); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3605 = 8'h8d == _T_24 ? $signed(regsA_71_im) : $signed(_GEN_3604); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3606 = 8'h8e == _T_24 ? $signed(regsA_72_im) : $signed(_GEN_3605); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3607 = 8'h8f == _T_24 ? $signed(regsA_73_im) : $signed(_GEN_3606); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3608 = 8'h90 == _T_24 ? $signed(regsA_74_im) : $signed(_GEN_3607); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3609 = 8'h91 == _T_24 ? $signed(regsA_75_im) : $signed(_GEN_3608); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3610 = 8'h92 == _T_24 ? $signed(regsA_76_im) : $signed(_GEN_3609); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3611 = 8'h93 == _T_24 ? $signed(regsA_77_im) : $signed(_GEN_3610); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3612 = 8'h94 == _T_24 ? $signed(regsA_78_im) : $signed(_GEN_3611); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3613 = 8'h95 == _T_24 ? $signed(regsA_79_im) : $signed(_GEN_3612); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3614 = 8'h96 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3613); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3615 = 8'h97 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3614); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3616 = 8'h98 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3615); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3617 = 8'h99 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3616); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3618 = 8'h9a == _T_24 ? $signed(32'sh0) : $signed(_GEN_3617); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3619 = 8'h9b == _T_24 ? $signed(32'sh0) : $signed(_GEN_3618); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3620 = 8'h9c == _T_24 ? $signed(32'sh0) : $signed(_GEN_3619); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3621 = 8'h9d == _T_24 ? $signed(32'sh0) : $signed(_GEN_3620); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3622 = 8'h9e == _T_24 ? $signed(32'sh0) : $signed(_GEN_3621); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3623 = 8'h9f == _T_24 ? $signed(32'sh0) : $signed(_GEN_3622); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3624 = 8'ha0 == _T_24 ? $signed(regsA_80_im) : $signed(_GEN_3623); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3625 = 8'ha1 == _T_24 ? $signed(regsA_81_im) : $signed(_GEN_3624); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3626 = 8'ha2 == _T_24 ? $signed(regsA_82_im) : $signed(_GEN_3625); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3627 = 8'ha3 == _T_24 ? $signed(regsA_83_im) : $signed(_GEN_3626); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3628 = 8'ha4 == _T_24 ? $signed(regsA_84_im) : $signed(_GEN_3627); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3629 = 8'ha5 == _T_24 ? $signed(regsA_85_im) : $signed(_GEN_3628); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3630 = 8'ha6 == _T_24 ? $signed(regsA_86_im) : $signed(_GEN_3629); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3631 = 8'ha7 == _T_24 ? $signed(regsA_87_im) : $signed(_GEN_3630); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3632 = 8'ha8 == _T_24 ? $signed(regsA_88_im) : $signed(_GEN_3631); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3633 = 8'ha9 == _T_24 ? $signed(regsA_89_im) : $signed(_GEN_3632); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3634 = 8'haa == _T_24 ? $signed(32'sh0) : $signed(_GEN_3633); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3635 = 8'hab == _T_24 ? $signed(32'sh0) : $signed(_GEN_3634); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3636 = 8'hac == _T_24 ? $signed(32'sh0) : $signed(_GEN_3635); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3637 = 8'had == _T_24 ? $signed(32'sh0) : $signed(_GEN_3636); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3638 = 8'hae == _T_24 ? $signed(32'sh0) : $signed(_GEN_3637); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3639 = 8'haf == _T_24 ? $signed(32'sh0) : $signed(_GEN_3638); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3640 = 8'hb0 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3639); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3641 = 8'hb1 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3640); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3642 = 8'hb2 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3641); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3643 = 8'hb3 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3642); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3644 = 8'hb4 == _T_24 ? $signed(regsA_90_im) : $signed(_GEN_3643); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3645 = 8'hb5 == _T_24 ? $signed(regsA_91_im) : $signed(_GEN_3644); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3646 = 8'hb6 == _T_24 ? $signed(regsA_92_im) : $signed(_GEN_3645); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3647 = 8'hb7 == _T_24 ? $signed(regsA_93_im) : $signed(_GEN_3646); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3648 = 8'hb8 == _T_24 ? $signed(regsA_94_im) : $signed(_GEN_3647); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3649 = 8'hb9 == _T_24 ? $signed(regsA_95_im) : $signed(_GEN_3648); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3650 = 8'hba == _T_24 ? $signed(regsA_96_im) : $signed(_GEN_3649); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3651 = 8'hbb == _T_24 ? $signed(regsA_97_im) : $signed(_GEN_3650); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3652 = 8'hbc == _T_24 ? $signed(regsA_98_im) : $signed(_GEN_3651); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3653 = 8'hbd == _T_24 ? $signed(regsA_99_im) : $signed(_GEN_3652); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3655 = 8'h1 == _T_24 ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3656 = 8'h2 == _T_24 ? $signed(regsA_2_re) : $signed(_GEN_3655); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3657 = 8'h3 == _T_24 ? $signed(regsA_3_re) : $signed(_GEN_3656); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3658 = 8'h4 == _T_24 ? $signed(regsA_4_re) : $signed(_GEN_3657); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3659 = 8'h5 == _T_24 ? $signed(regsA_5_re) : $signed(_GEN_3658); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3660 = 8'h6 == _T_24 ? $signed(regsA_6_re) : $signed(_GEN_3659); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3661 = 8'h7 == _T_24 ? $signed(regsA_7_re) : $signed(_GEN_3660); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3662 = 8'h8 == _T_24 ? $signed(regsA_8_re) : $signed(_GEN_3661); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3663 = 8'h9 == _T_24 ? $signed(regsA_9_re) : $signed(_GEN_3662); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3664 = 8'ha == _T_24 ? $signed(32'sh0) : $signed(_GEN_3663); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3665 = 8'hb == _T_24 ? $signed(32'sh0) : $signed(_GEN_3664); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3666 = 8'hc == _T_24 ? $signed(32'sh0) : $signed(_GEN_3665); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3667 = 8'hd == _T_24 ? $signed(32'sh0) : $signed(_GEN_3666); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3668 = 8'he == _T_24 ? $signed(32'sh0) : $signed(_GEN_3667); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3669 = 8'hf == _T_24 ? $signed(32'sh0) : $signed(_GEN_3668); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3670 = 8'h10 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3669); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3671 = 8'h11 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3670); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3672 = 8'h12 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3671); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3673 = 8'h13 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3672); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3674 = 8'h14 == _T_24 ? $signed(regsA_10_re) : $signed(_GEN_3673); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3675 = 8'h15 == _T_24 ? $signed(regsA_11_re) : $signed(_GEN_3674); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3676 = 8'h16 == _T_24 ? $signed(regsA_12_re) : $signed(_GEN_3675); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3677 = 8'h17 == _T_24 ? $signed(regsA_13_re) : $signed(_GEN_3676); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3678 = 8'h18 == _T_24 ? $signed(regsA_14_re) : $signed(_GEN_3677); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3679 = 8'h19 == _T_24 ? $signed(regsA_15_re) : $signed(_GEN_3678); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3680 = 8'h1a == _T_24 ? $signed(regsA_16_re) : $signed(_GEN_3679); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3681 = 8'h1b == _T_24 ? $signed(regsA_17_re) : $signed(_GEN_3680); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3682 = 8'h1c == _T_24 ? $signed(regsA_18_re) : $signed(_GEN_3681); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3683 = 8'h1d == _T_24 ? $signed(regsA_19_re) : $signed(_GEN_3682); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3684 = 8'h1e == _T_24 ? $signed(32'sh0) : $signed(_GEN_3683); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3685 = 8'h1f == _T_24 ? $signed(32'sh0) : $signed(_GEN_3684); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3686 = 8'h20 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3685); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3687 = 8'h21 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3686); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3688 = 8'h22 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3687); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3689 = 8'h23 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3688); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3690 = 8'h24 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3689); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3691 = 8'h25 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3690); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3692 = 8'h26 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3691); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3693 = 8'h27 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3692); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3694 = 8'h28 == _T_24 ? $signed(regsA_20_re) : $signed(_GEN_3693); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3695 = 8'h29 == _T_24 ? $signed(regsA_21_re) : $signed(_GEN_3694); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3696 = 8'h2a == _T_24 ? $signed(regsA_22_re) : $signed(_GEN_3695); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3697 = 8'h2b == _T_24 ? $signed(regsA_23_re) : $signed(_GEN_3696); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3698 = 8'h2c == _T_24 ? $signed(regsA_24_re) : $signed(_GEN_3697); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3699 = 8'h2d == _T_24 ? $signed(regsA_25_re) : $signed(_GEN_3698); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3700 = 8'h2e == _T_24 ? $signed(regsA_26_re) : $signed(_GEN_3699); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3701 = 8'h2f == _T_24 ? $signed(regsA_27_re) : $signed(_GEN_3700); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3702 = 8'h30 == _T_24 ? $signed(regsA_28_re) : $signed(_GEN_3701); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3703 = 8'h31 == _T_24 ? $signed(regsA_29_re) : $signed(_GEN_3702); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3704 = 8'h32 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3703); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3705 = 8'h33 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3704); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3706 = 8'h34 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3705); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3707 = 8'h35 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3706); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3708 = 8'h36 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3707); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3709 = 8'h37 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3708); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3710 = 8'h38 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3709); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3711 = 8'h39 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3710); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3712 = 8'h3a == _T_24 ? $signed(32'sh0) : $signed(_GEN_3711); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3713 = 8'h3b == _T_24 ? $signed(32'sh0) : $signed(_GEN_3712); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3714 = 8'h3c == _T_24 ? $signed(regsA_30_re) : $signed(_GEN_3713); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3715 = 8'h3d == _T_24 ? $signed(regsA_31_re) : $signed(_GEN_3714); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3716 = 8'h3e == _T_24 ? $signed(regsA_32_re) : $signed(_GEN_3715); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3717 = 8'h3f == _T_24 ? $signed(regsA_33_re) : $signed(_GEN_3716); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3718 = 8'h40 == _T_24 ? $signed(regsA_34_re) : $signed(_GEN_3717); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3719 = 8'h41 == _T_24 ? $signed(regsA_35_re) : $signed(_GEN_3718); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3720 = 8'h42 == _T_24 ? $signed(regsA_36_re) : $signed(_GEN_3719); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3721 = 8'h43 == _T_24 ? $signed(regsA_37_re) : $signed(_GEN_3720); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3722 = 8'h44 == _T_24 ? $signed(regsA_38_re) : $signed(_GEN_3721); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3723 = 8'h45 == _T_24 ? $signed(regsA_39_re) : $signed(_GEN_3722); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3724 = 8'h46 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3723); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3725 = 8'h47 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3724); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3726 = 8'h48 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3725); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3727 = 8'h49 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3726); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3728 = 8'h4a == _T_24 ? $signed(32'sh0) : $signed(_GEN_3727); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3729 = 8'h4b == _T_24 ? $signed(32'sh0) : $signed(_GEN_3728); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3730 = 8'h4c == _T_24 ? $signed(32'sh0) : $signed(_GEN_3729); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3731 = 8'h4d == _T_24 ? $signed(32'sh0) : $signed(_GEN_3730); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3732 = 8'h4e == _T_24 ? $signed(32'sh0) : $signed(_GEN_3731); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3733 = 8'h4f == _T_24 ? $signed(32'sh0) : $signed(_GEN_3732); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3734 = 8'h50 == _T_24 ? $signed(regsA_40_re) : $signed(_GEN_3733); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3735 = 8'h51 == _T_24 ? $signed(regsA_41_re) : $signed(_GEN_3734); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3736 = 8'h52 == _T_24 ? $signed(regsA_42_re) : $signed(_GEN_3735); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3737 = 8'h53 == _T_24 ? $signed(regsA_43_re) : $signed(_GEN_3736); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3738 = 8'h54 == _T_24 ? $signed(regsA_44_re) : $signed(_GEN_3737); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3739 = 8'h55 == _T_24 ? $signed(regsA_45_re) : $signed(_GEN_3738); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3740 = 8'h56 == _T_24 ? $signed(regsA_46_re) : $signed(_GEN_3739); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3741 = 8'h57 == _T_24 ? $signed(regsA_47_re) : $signed(_GEN_3740); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3742 = 8'h58 == _T_24 ? $signed(regsA_48_re) : $signed(_GEN_3741); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3743 = 8'h59 == _T_24 ? $signed(regsA_49_re) : $signed(_GEN_3742); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3744 = 8'h5a == _T_24 ? $signed(32'sh0) : $signed(_GEN_3743); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3745 = 8'h5b == _T_24 ? $signed(32'sh0) : $signed(_GEN_3744); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3746 = 8'h5c == _T_24 ? $signed(32'sh0) : $signed(_GEN_3745); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3747 = 8'h5d == _T_24 ? $signed(32'sh0) : $signed(_GEN_3746); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3748 = 8'h5e == _T_24 ? $signed(32'sh0) : $signed(_GEN_3747); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3749 = 8'h5f == _T_24 ? $signed(32'sh0) : $signed(_GEN_3748); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3750 = 8'h60 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3749); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3751 = 8'h61 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3750); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3752 = 8'h62 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3751); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3753 = 8'h63 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3752); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3754 = 8'h64 == _T_24 ? $signed(regsA_50_re) : $signed(_GEN_3753); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3755 = 8'h65 == _T_24 ? $signed(regsA_51_re) : $signed(_GEN_3754); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3756 = 8'h66 == _T_24 ? $signed(regsA_52_re) : $signed(_GEN_3755); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3757 = 8'h67 == _T_24 ? $signed(regsA_53_re) : $signed(_GEN_3756); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3758 = 8'h68 == _T_24 ? $signed(regsA_54_re) : $signed(_GEN_3757); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3759 = 8'h69 == _T_24 ? $signed(regsA_55_re) : $signed(_GEN_3758); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3760 = 8'h6a == _T_24 ? $signed(regsA_56_re) : $signed(_GEN_3759); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3761 = 8'h6b == _T_24 ? $signed(regsA_57_re) : $signed(_GEN_3760); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3762 = 8'h6c == _T_24 ? $signed(regsA_58_re) : $signed(_GEN_3761); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3763 = 8'h6d == _T_24 ? $signed(regsA_59_re) : $signed(_GEN_3762); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3764 = 8'h6e == _T_24 ? $signed(32'sh0) : $signed(_GEN_3763); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3765 = 8'h6f == _T_24 ? $signed(32'sh0) : $signed(_GEN_3764); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3766 = 8'h70 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3765); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3767 = 8'h71 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3766); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3768 = 8'h72 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3767); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3769 = 8'h73 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3768); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3770 = 8'h74 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3769); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3771 = 8'h75 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3770); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3772 = 8'h76 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3771); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3773 = 8'h77 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3772); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3774 = 8'h78 == _T_24 ? $signed(regsA_60_re) : $signed(_GEN_3773); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3775 = 8'h79 == _T_24 ? $signed(regsA_61_re) : $signed(_GEN_3774); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3776 = 8'h7a == _T_24 ? $signed(regsA_62_re) : $signed(_GEN_3775); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3777 = 8'h7b == _T_24 ? $signed(regsA_63_re) : $signed(_GEN_3776); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3778 = 8'h7c == _T_24 ? $signed(regsA_64_re) : $signed(_GEN_3777); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3779 = 8'h7d == _T_24 ? $signed(regsA_65_re) : $signed(_GEN_3778); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3780 = 8'h7e == _T_24 ? $signed(regsA_66_re) : $signed(_GEN_3779); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3781 = 8'h7f == _T_24 ? $signed(regsA_67_re) : $signed(_GEN_3780); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3782 = 8'h80 == _T_24 ? $signed(regsA_68_re) : $signed(_GEN_3781); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3783 = 8'h81 == _T_24 ? $signed(regsA_69_re) : $signed(_GEN_3782); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3784 = 8'h82 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3783); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3785 = 8'h83 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3784); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3786 = 8'h84 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3785); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3787 = 8'h85 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3786); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3788 = 8'h86 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3787); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3789 = 8'h87 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3788); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3790 = 8'h88 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3789); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3791 = 8'h89 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3790); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3792 = 8'h8a == _T_24 ? $signed(32'sh0) : $signed(_GEN_3791); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3793 = 8'h8b == _T_24 ? $signed(32'sh0) : $signed(_GEN_3792); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3794 = 8'h8c == _T_24 ? $signed(regsA_70_re) : $signed(_GEN_3793); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3795 = 8'h8d == _T_24 ? $signed(regsA_71_re) : $signed(_GEN_3794); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3796 = 8'h8e == _T_24 ? $signed(regsA_72_re) : $signed(_GEN_3795); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3797 = 8'h8f == _T_24 ? $signed(regsA_73_re) : $signed(_GEN_3796); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3798 = 8'h90 == _T_24 ? $signed(regsA_74_re) : $signed(_GEN_3797); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3799 = 8'h91 == _T_24 ? $signed(regsA_75_re) : $signed(_GEN_3798); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3800 = 8'h92 == _T_24 ? $signed(regsA_76_re) : $signed(_GEN_3799); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3801 = 8'h93 == _T_24 ? $signed(regsA_77_re) : $signed(_GEN_3800); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3802 = 8'h94 == _T_24 ? $signed(regsA_78_re) : $signed(_GEN_3801); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3803 = 8'h95 == _T_24 ? $signed(regsA_79_re) : $signed(_GEN_3802); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3804 = 8'h96 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3803); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3805 = 8'h97 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3804); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3806 = 8'h98 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3805); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3807 = 8'h99 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3806); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3808 = 8'h9a == _T_24 ? $signed(32'sh0) : $signed(_GEN_3807); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3809 = 8'h9b == _T_24 ? $signed(32'sh0) : $signed(_GEN_3808); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3810 = 8'h9c == _T_24 ? $signed(32'sh0) : $signed(_GEN_3809); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3811 = 8'h9d == _T_24 ? $signed(32'sh0) : $signed(_GEN_3810); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3812 = 8'h9e == _T_24 ? $signed(32'sh0) : $signed(_GEN_3811); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3813 = 8'h9f == _T_24 ? $signed(32'sh0) : $signed(_GEN_3812); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3814 = 8'ha0 == _T_24 ? $signed(regsA_80_re) : $signed(_GEN_3813); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3815 = 8'ha1 == _T_24 ? $signed(regsA_81_re) : $signed(_GEN_3814); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3816 = 8'ha2 == _T_24 ? $signed(regsA_82_re) : $signed(_GEN_3815); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3817 = 8'ha3 == _T_24 ? $signed(regsA_83_re) : $signed(_GEN_3816); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3818 = 8'ha4 == _T_24 ? $signed(regsA_84_re) : $signed(_GEN_3817); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3819 = 8'ha5 == _T_24 ? $signed(regsA_85_re) : $signed(_GEN_3818); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3820 = 8'ha6 == _T_24 ? $signed(regsA_86_re) : $signed(_GEN_3819); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3821 = 8'ha7 == _T_24 ? $signed(regsA_87_re) : $signed(_GEN_3820); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3822 = 8'ha8 == _T_24 ? $signed(regsA_88_re) : $signed(_GEN_3821); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3823 = 8'ha9 == _T_24 ? $signed(regsA_89_re) : $signed(_GEN_3822); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3824 = 8'haa == _T_24 ? $signed(32'sh0) : $signed(_GEN_3823); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3825 = 8'hab == _T_24 ? $signed(32'sh0) : $signed(_GEN_3824); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3826 = 8'hac == _T_24 ? $signed(32'sh0) : $signed(_GEN_3825); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3827 = 8'had == _T_24 ? $signed(32'sh0) : $signed(_GEN_3826); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3828 = 8'hae == _T_24 ? $signed(32'sh0) : $signed(_GEN_3827); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3829 = 8'haf == _T_24 ? $signed(32'sh0) : $signed(_GEN_3828); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3830 = 8'hb0 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3829); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3831 = 8'hb1 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3830); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3832 = 8'hb2 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3831); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3833 = 8'hb3 == _T_24 ? $signed(32'sh0) : $signed(_GEN_3832); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3834 = 8'hb4 == _T_24 ? $signed(regsA_90_re) : $signed(_GEN_3833); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3835 = 8'hb5 == _T_24 ? $signed(regsA_91_re) : $signed(_GEN_3834); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3836 = 8'hb6 == _T_24 ? $signed(regsA_92_re) : $signed(_GEN_3835); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3837 = 8'hb7 == _T_24 ? $signed(regsA_93_re) : $signed(_GEN_3836); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3838 = 8'hb8 == _T_24 ? $signed(regsA_94_re) : $signed(_GEN_3837); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3839 = 8'hb9 == _T_24 ? $signed(regsA_95_re) : $signed(_GEN_3838); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3840 = 8'hba == _T_24 ? $signed(regsA_96_re) : $signed(_GEN_3839); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3841 = 8'hbb == _T_24 ? $signed(regsA_97_re) : $signed(_GEN_3840); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3842 = 8'hbc == _T_24 ? $signed(regsA_98_re) : $signed(_GEN_3841); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3843 = 8'hbd == _T_24 ? $signed(regsA_99_re) : $signed(_GEN_3842); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [8:0] _T_25 = 4'h8 * 5'h13; // @[Matrix_Mul_V1.scala 148:44]
  wire [8:0] _GEN_9203 = {{3'd0}, input_point}; // @[Matrix_Mul_V1.scala 148:60]
  wire [8:0] _T_27 = _T_25 + _GEN_9203; // @[Matrix_Mul_V1.scala 148:60]
  wire [31:0] _GEN_3845 = 8'h1 == _T_27[7:0] ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3846 = 8'h2 == _T_27[7:0] ? $signed(regsA_2_im) : $signed(_GEN_3845); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3847 = 8'h3 == _T_27[7:0] ? $signed(regsA_3_im) : $signed(_GEN_3846); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3848 = 8'h4 == _T_27[7:0] ? $signed(regsA_4_im) : $signed(_GEN_3847); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3849 = 8'h5 == _T_27[7:0] ? $signed(regsA_5_im) : $signed(_GEN_3848); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3850 = 8'h6 == _T_27[7:0] ? $signed(regsA_6_im) : $signed(_GEN_3849); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3851 = 8'h7 == _T_27[7:0] ? $signed(regsA_7_im) : $signed(_GEN_3850); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3852 = 8'h8 == _T_27[7:0] ? $signed(regsA_8_im) : $signed(_GEN_3851); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3853 = 8'h9 == _T_27[7:0] ? $signed(regsA_9_im) : $signed(_GEN_3852); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3854 = 8'ha == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3853); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3855 = 8'hb == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3854); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3856 = 8'hc == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3855); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3857 = 8'hd == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3856); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3858 = 8'he == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3857); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3859 = 8'hf == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3858); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3860 = 8'h10 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3859); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3861 = 8'h11 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3860); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3862 = 8'h12 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3861); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3863 = 8'h13 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3862); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3864 = 8'h14 == _T_27[7:0] ? $signed(regsA_10_im) : $signed(_GEN_3863); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3865 = 8'h15 == _T_27[7:0] ? $signed(regsA_11_im) : $signed(_GEN_3864); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3866 = 8'h16 == _T_27[7:0] ? $signed(regsA_12_im) : $signed(_GEN_3865); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3867 = 8'h17 == _T_27[7:0] ? $signed(regsA_13_im) : $signed(_GEN_3866); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3868 = 8'h18 == _T_27[7:0] ? $signed(regsA_14_im) : $signed(_GEN_3867); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3869 = 8'h19 == _T_27[7:0] ? $signed(regsA_15_im) : $signed(_GEN_3868); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3870 = 8'h1a == _T_27[7:0] ? $signed(regsA_16_im) : $signed(_GEN_3869); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3871 = 8'h1b == _T_27[7:0] ? $signed(regsA_17_im) : $signed(_GEN_3870); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3872 = 8'h1c == _T_27[7:0] ? $signed(regsA_18_im) : $signed(_GEN_3871); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3873 = 8'h1d == _T_27[7:0] ? $signed(regsA_19_im) : $signed(_GEN_3872); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3874 = 8'h1e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3873); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3875 = 8'h1f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3874); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3876 = 8'h20 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3875); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3877 = 8'h21 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3876); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3878 = 8'h22 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3877); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3879 = 8'h23 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3878); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3880 = 8'h24 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3879); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3881 = 8'h25 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3880); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3882 = 8'h26 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3881); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3883 = 8'h27 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3882); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3884 = 8'h28 == _T_27[7:0] ? $signed(regsA_20_im) : $signed(_GEN_3883); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3885 = 8'h29 == _T_27[7:0] ? $signed(regsA_21_im) : $signed(_GEN_3884); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3886 = 8'h2a == _T_27[7:0] ? $signed(regsA_22_im) : $signed(_GEN_3885); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3887 = 8'h2b == _T_27[7:0] ? $signed(regsA_23_im) : $signed(_GEN_3886); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3888 = 8'h2c == _T_27[7:0] ? $signed(regsA_24_im) : $signed(_GEN_3887); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3889 = 8'h2d == _T_27[7:0] ? $signed(regsA_25_im) : $signed(_GEN_3888); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3890 = 8'h2e == _T_27[7:0] ? $signed(regsA_26_im) : $signed(_GEN_3889); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3891 = 8'h2f == _T_27[7:0] ? $signed(regsA_27_im) : $signed(_GEN_3890); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3892 = 8'h30 == _T_27[7:0] ? $signed(regsA_28_im) : $signed(_GEN_3891); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3893 = 8'h31 == _T_27[7:0] ? $signed(regsA_29_im) : $signed(_GEN_3892); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3894 = 8'h32 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3893); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3895 = 8'h33 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3894); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3896 = 8'h34 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3895); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3897 = 8'h35 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3896); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3898 = 8'h36 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3897); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3899 = 8'h37 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3898); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3900 = 8'h38 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3899); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3901 = 8'h39 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3900); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3902 = 8'h3a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3901); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3903 = 8'h3b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3902); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3904 = 8'h3c == _T_27[7:0] ? $signed(regsA_30_im) : $signed(_GEN_3903); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3905 = 8'h3d == _T_27[7:0] ? $signed(regsA_31_im) : $signed(_GEN_3904); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3906 = 8'h3e == _T_27[7:0] ? $signed(regsA_32_im) : $signed(_GEN_3905); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3907 = 8'h3f == _T_27[7:0] ? $signed(regsA_33_im) : $signed(_GEN_3906); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3908 = 8'h40 == _T_27[7:0] ? $signed(regsA_34_im) : $signed(_GEN_3907); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3909 = 8'h41 == _T_27[7:0] ? $signed(regsA_35_im) : $signed(_GEN_3908); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3910 = 8'h42 == _T_27[7:0] ? $signed(regsA_36_im) : $signed(_GEN_3909); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3911 = 8'h43 == _T_27[7:0] ? $signed(regsA_37_im) : $signed(_GEN_3910); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3912 = 8'h44 == _T_27[7:0] ? $signed(regsA_38_im) : $signed(_GEN_3911); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3913 = 8'h45 == _T_27[7:0] ? $signed(regsA_39_im) : $signed(_GEN_3912); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3914 = 8'h46 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3913); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3915 = 8'h47 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3914); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3916 = 8'h48 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3915); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3917 = 8'h49 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3916); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3918 = 8'h4a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3917); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3919 = 8'h4b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3918); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3920 = 8'h4c == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3919); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3921 = 8'h4d == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3920); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3922 = 8'h4e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3921); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3923 = 8'h4f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3922); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3924 = 8'h50 == _T_27[7:0] ? $signed(regsA_40_im) : $signed(_GEN_3923); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3925 = 8'h51 == _T_27[7:0] ? $signed(regsA_41_im) : $signed(_GEN_3924); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3926 = 8'h52 == _T_27[7:0] ? $signed(regsA_42_im) : $signed(_GEN_3925); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3927 = 8'h53 == _T_27[7:0] ? $signed(regsA_43_im) : $signed(_GEN_3926); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3928 = 8'h54 == _T_27[7:0] ? $signed(regsA_44_im) : $signed(_GEN_3927); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3929 = 8'h55 == _T_27[7:0] ? $signed(regsA_45_im) : $signed(_GEN_3928); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3930 = 8'h56 == _T_27[7:0] ? $signed(regsA_46_im) : $signed(_GEN_3929); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3931 = 8'h57 == _T_27[7:0] ? $signed(regsA_47_im) : $signed(_GEN_3930); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3932 = 8'h58 == _T_27[7:0] ? $signed(regsA_48_im) : $signed(_GEN_3931); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3933 = 8'h59 == _T_27[7:0] ? $signed(regsA_49_im) : $signed(_GEN_3932); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3934 = 8'h5a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3933); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3935 = 8'h5b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3934); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3936 = 8'h5c == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3935); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3937 = 8'h5d == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3936); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3938 = 8'h5e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3937); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3939 = 8'h5f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3938); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3940 = 8'h60 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3939); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3941 = 8'h61 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3940); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3942 = 8'h62 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3941); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3943 = 8'h63 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3942); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3944 = 8'h64 == _T_27[7:0] ? $signed(regsA_50_im) : $signed(_GEN_3943); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3945 = 8'h65 == _T_27[7:0] ? $signed(regsA_51_im) : $signed(_GEN_3944); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3946 = 8'h66 == _T_27[7:0] ? $signed(regsA_52_im) : $signed(_GEN_3945); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3947 = 8'h67 == _T_27[7:0] ? $signed(regsA_53_im) : $signed(_GEN_3946); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3948 = 8'h68 == _T_27[7:0] ? $signed(regsA_54_im) : $signed(_GEN_3947); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3949 = 8'h69 == _T_27[7:0] ? $signed(regsA_55_im) : $signed(_GEN_3948); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3950 = 8'h6a == _T_27[7:0] ? $signed(regsA_56_im) : $signed(_GEN_3949); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3951 = 8'h6b == _T_27[7:0] ? $signed(regsA_57_im) : $signed(_GEN_3950); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3952 = 8'h6c == _T_27[7:0] ? $signed(regsA_58_im) : $signed(_GEN_3951); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3953 = 8'h6d == _T_27[7:0] ? $signed(regsA_59_im) : $signed(_GEN_3952); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3954 = 8'h6e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3953); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3955 = 8'h6f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3954); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3956 = 8'h70 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3955); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3957 = 8'h71 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3956); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3958 = 8'h72 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3957); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3959 = 8'h73 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3958); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3960 = 8'h74 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3959); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3961 = 8'h75 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3960); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3962 = 8'h76 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3961); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3963 = 8'h77 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3962); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3964 = 8'h78 == _T_27[7:0] ? $signed(regsA_60_im) : $signed(_GEN_3963); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3965 = 8'h79 == _T_27[7:0] ? $signed(regsA_61_im) : $signed(_GEN_3964); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3966 = 8'h7a == _T_27[7:0] ? $signed(regsA_62_im) : $signed(_GEN_3965); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3967 = 8'h7b == _T_27[7:0] ? $signed(regsA_63_im) : $signed(_GEN_3966); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3968 = 8'h7c == _T_27[7:0] ? $signed(regsA_64_im) : $signed(_GEN_3967); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3969 = 8'h7d == _T_27[7:0] ? $signed(regsA_65_im) : $signed(_GEN_3968); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3970 = 8'h7e == _T_27[7:0] ? $signed(regsA_66_im) : $signed(_GEN_3969); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3971 = 8'h7f == _T_27[7:0] ? $signed(regsA_67_im) : $signed(_GEN_3970); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3972 = 8'h80 == _T_27[7:0] ? $signed(regsA_68_im) : $signed(_GEN_3971); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3973 = 8'h81 == _T_27[7:0] ? $signed(regsA_69_im) : $signed(_GEN_3972); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3974 = 8'h82 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3973); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3975 = 8'h83 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3974); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3976 = 8'h84 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3975); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3977 = 8'h85 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3976); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3978 = 8'h86 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3977); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3979 = 8'h87 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3978); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3980 = 8'h88 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3979); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3981 = 8'h89 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3980); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3982 = 8'h8a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3981); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3983 = 8'h8b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3982); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3984 = 8'h8c == _T_27[7:0] ? $signed(regsA_70_im) : $signed(_GEN_3983); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3985 = 8'h8d == _T_27[7:0] ? $signed(regsA_71_im) : $signed(_GEN_3984); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3986 = 8'h8e == _T_27[7:0] ? $signed(regsA_72_im) : $signed(_GEN_3985); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3987 = 8'h8f == _T_27[7:0] ? $signed(regsA_73_im) : $signed(_GEN_3986); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3988 = 8'h90 == _T_27[7:0] ? $signed(regsA_74_im) : $signed(_GEN_3987); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3989 = 8'h91 == _T_27[7:0] ? $signed(regsA_75_im) : $signed(_GEN_3988); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3990 = 8'h92 == _T_27[7:0] ? $signed(regsA_76_im) : $signed(_GEN_3989); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3991 = 8'h93 == _T_27[7:0] ? $signed(regsA_77_im) : $signed(_GEN_3990); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3992 = 8'h94 == _T_27[7:0] ? $signed(regsA_78_im) : $signed(_GEN_3991); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3993 = 8'h95 == _T_27[7:0] ? $signed(regsA_79_im) : $signed(_GEN_3992); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3994 = 8'h96 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3993); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3995 = 8'h97 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3994); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3996 = 8'h98 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3995); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3997 = 8'h99 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3996); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3998 = 8'h9a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3997); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_3999 = 8'h9b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3998); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4000 = 8'h9c == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_3999); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4001 = 8'h9d == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4000); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4002 = 8'h9e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4001); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4003 = 8'h9f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4002); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4004 = 8'ha0 == _T_27[7:0] ? $signed(regsA_80_im) : $signed(_GEN_4003); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4005 = 8'ha1 == _T_27[7:0] ? $signed(regsA_81_im) : $signed(_GEN_4004); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4006 = 8'ha2 == _T_27[7:0] ? $signed(regsA_82_im) : $signed(_GEN_4005); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4007 = 8'ha3 == _T_27[7:0] ? $signed(regsA_83_im) : $signed(_GEN_4006); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4008 = 8'ha4 == _T_27[7:0] ? $signed(regsA_84_im) : $signed(_GEN_4007); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4009 = 8'ha5 == _T_27[7:0] ? $signed(regsA_85_im) : $signed(_GEN_4008); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4010 = 8'ha6 == _T_27[7:0] ? $signed(regsA_86_im) : $signed(_GEN_4009); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4011 = 8'ha7 == _T_27[7:0] ? $signed(regsA_87_im) : $signed(_GEN_4010); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4012 = 8'ha8 == _T_27[7:0] ? $signed(regsA_88_im) : $signed(_GEN_4011); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4013 = 8'ha9 == _T_27[7:0] ? $signed(regsA_89_im) : $signed(_GEN_4012); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4014 = 8'haa == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4013); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4015 = 8'hab == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4014); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4016 = 8'hac == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4015); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4017 = 8'had == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4016); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4018 = 8'hae == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4017); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4019 = 8'haf == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4018); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4020 = 8'hb0 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4019); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4021 = 8'hb1 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4020); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4022 = 8'hb2 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4021); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4023 = 8'hb3 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4022); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4024 = 8'hb4 == _T_27[7:0] ? $signed(regsA_90_im) : $signed(_GEN_4023); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4025 = 8'hb5 == _T_27[7:0] ? $signed(regsA_91_im) : $signed(_GEN_4024); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4026 = 8'hb6 == _T_27[7:0] ? $signed(regsA_92_im) : $signed(_GEN_4025); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4027 = 8'hb7 == _T_27[7:0] ? $signed(regsA_93_im) : $signed(_GEN_4026); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4028 = 8'hb8 == _T_27[7:0] ? $signed(regsA_94_im) : $signed(_GEN_4027); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4029 = 8'hb9 == _T_27[7:0] ? $signed(regsA_95_im) : $signed(_GEN_4028); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4030 = 8'hba == _T_27[7:0] ? $signed(regsA_96_im) : $signed(_GEN_4029); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4031 = 8'hbb == _T_27[7:0] ? $signed(regsA_97_im) : $signed(_GEN_4030); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4032 = 8'hbc == _T_27[7:0] ? $signed(regsA_98_im) : $signed(_GEN_4031); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4033 = 8'hbd == _T_27[7:0] ? $signed(regsA_99_im) : $signed(_GEN_4032); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4035 = 8'h1 == _T_27[7:0] ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4036 = 8'h2 == _T_27[7:0] ? $signed(regsA_2_re) : $signed(_GEN_4035); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4037 = 8'h3 == _T_27[7:0] ? $signed(regsA_3_re) : $signed(_GEN_4036); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4038 = 8'h4 == _T_27[7:0] ? $signed(regsA_4_re) : $signed(_GEN_4037); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4039 = 8'h5 == _T_27[7:0] ? $signed(regsA_5_re) : $signed(_GEN_4038); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4040 = 8'h6 == _T_27[7:0] ? $signed(regsA_6_re) : $signed(_GEN_4039); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4041 = 8'h7 == _T_27[7:0] ? $signed(regsA_7_re) : $signed(_GEN_4040); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4042 = 8'h8 == _T_27[7:0] ? $signed(regsA_8_re) : $signed(_GEN_4041); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4043 = 8'h9 == _T_27[7:0] ? $signed(regsA_9_re) : $signed(_GEN_4042); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4044 = 8'ha == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4043); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4045 = 8'hb == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4044); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4046 = 8'hc == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4045); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4047 = 8'hd == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4046); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4048 = 8'he == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4047); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4049 = 8'hf == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4048); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4050 = 8'h10 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4049); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4051 = 8'h11 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4050); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4052 = 8'h12 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4051); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4053 = 8'h13 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4052); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4054 = 8'h14 == _T_27[7:0] ? $signed(regsA_10_re) : $signed(_GEN_4053); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4055 = 8'h15 == _T_27[7:0] ? $signed(regsA_11_re) : $signed(_GEN_4054); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4056 = 8'h16 == _T_27[7:0] ? $signed(regsA_12_re) : $signed(_GEN_4055); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4057 = 8'h17 == _T_27[7:0] ? $signed(regsA_13_re) : $signed(_GEN_4056); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4058 = 8'h18 == _T_27[7:0] ? $signed(regsA_14_re) : $signed(_GEN_4057); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4059 = 8'h19 == _T_27[7:0] ? $signed(regsA_15_re) : $signed(_GEN_4058); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4060 = 8'h1a == _T_27[7:0] ? $signed(regsA_16_re) : $signed(_GEN_4059); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4061 = 8'h1b == _T_27[7:0] ? $signed(regsA_17_re) : $signed(_GEN_4060); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4062 = 8'h1c == _T_27[7:0] ? $signed(regsA_18_re) : $signed(_GEN_4061); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4063 = 8'h1d == _T_27[7:0] ? $signed(regsA_19_re) : $signed(_GEN_4062); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4064 = 8'h1e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4063); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4065 = 8'h1f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4064); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4066 = 8'h20 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4065); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4067 = 8'h21 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4066); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4068 = 8'h22 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4067); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4069 = 8'h23 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4068); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4070 = 8'h24 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4069); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4071 = 8'h25 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4070); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4072 = 8'h26 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4071); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4073 = 8'h27 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4072); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4074 = 8'h28 == _T_27[7:0] ? $signed(regsA_20_re) : $signed(_GEN_4073); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4075 = 8'h29 == _T_27[7:0] ? $signed(regsA_21_re) : $signed(_GEN_4074); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4076 = 8'h2a == _T_27[7:0] ? $signed(regsA_22_re) : $signed(_GEN_4075); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4077 = 8'h2b == _T_27[7:0] ? $signed(regsA_23_re) : $signed(_GEN_4076); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4078 = 8'h2c == _T_27[7:0] ? $signed(regsA_24_re) : $signed(_GEN_4077); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4079 = 8'h2d == _T_27[7:0] ? $signed(regsA_25_re) : $signed(_GEN_4078); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4080 = 8'h2e == _T_27[7:0] ? $signed(regsA_26_re) : $signed(_GEN_4079); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4081 = 8'h2f == _T_27[7:0] ? $signed(regsA_27_re) : $signed(_GEN_4080); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4082 = 8'h30 == _T_27[7:0] ? $signed(regsA_28_re) : $signed(_GEN_4081); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4083 = 8'h31 == _T_27[7:0] ? $signed(regsA_29_re) : $signed(_GEN_4082); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4084 = 8'h32 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4083); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4085 = 8'h33 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4084); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4086 = 8'h34 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4085); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4087 = 8'h35 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4086); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4088 = 8'h36 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4087); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4089 = 8'h37 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4088); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4090 = 8'h38 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4089); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4091 = 8'h39 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4090); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4092 = 8'h3a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4091); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4093 = 8'h3b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4092); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4094 = 8'h3c == _T_27[7:0] ? $signed(regsA_30_re) : $signed(_GEN_4093); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4095 = 8'h3d == _T_27[7:0] ? $signed(regsA_31_re) : $signed(_GEN_4094); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4096 = 8'h3e == _T_27[7:0] ? $signed(regsA_32_re) : $signed(_GEN_4095); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4097 = 8'h3f == _T_27[7:0] ? $signed(regsA_33_re) : $signed(_GEN_4096); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4098 = 8'h40 == _T_27[7:0] ? $signed(regsA_34_re) : $signed(_GEN_4097); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4099 = 8'h41 == _T_27[7:0] ? $signed(regsA_35_re) : $signed(_GEN_4098); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4100 = 8'h42 == _T_27[7:0] ? $signed(regsA_36_re) : $signed(_GEN_4099); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4101 = 8'h43 == _T_27[7:0] ? $signed(regsA_37_re) : $signed(_GEN_4100); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4102 = 8'h44 == _T_27[7:0] ? $signed(regsA_38_re) : $signed(_GEN_4101); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4103 = 8'h45 == _T_27[7:0] ? $signed(regsA_39_re) : $signed(_GEN_4102); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4104 = 8'h46 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4103); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4105 = 8'h47 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4104); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4106 = 8'h48 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4105); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4107 = 8'h49 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4106); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4108 = 8'h4a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4107); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4109 = 8'h4b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4108); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4110 = 8'h4c == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4109); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4111 = 8'h4d == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4110); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4112 = 8'h4e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4111); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4113 = 8'h4f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4112); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4114 = 8'h50 == _T_27[7:0] ? $signed(regsA_40_re) : $signed(_GEN_4113); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4115 = 8'h51 == _T_27[7:0] ? $signed(regsA_41_re) : $signed(_GEN_4114); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4116 = 8'h52 == _T_27[7:0] ? $signed(regsA_42_re) : $signed(_GEN_4115); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4117 = 8'h53 == _T_27[7:0] ? $signed(regsA_43_re) : $signed(_GEN_4116); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4118 = 8'h54 == _T_27[7:0] ? $signed(regsA_44_re) : $signed(_GEN_4117); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4119 = 8'h55 == _T_27[7:0] ? $signed(regsA_45_re) : $signed(_GEN_4118); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4120 = 8'h56 == _T_27[7:0] ? $signed(regsA_46_re) : $signed(_GEN_4119); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4121 = 8'h57 == _T_27[7:0] ? $signed(regsA_47_re) : $signed(_GEN_4120); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4122 = 8'h58 == _T_27[7:0] ? $signed(regsA_48_re) : $signed(_GEN_4121); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4123 = 8'h59 == _T_27[7:0] ? $signed(regsA_49_re) : $signed(_GEN_4122); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4124 = 8'h5a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4123); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4125 = 8'h5b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4124); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4126 = 8'h5c == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4125); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4127 = 8'h5d == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4126); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4128 = 8'h5e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4127); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4129 = 8'h5f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4128); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4130 = 8'h60 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4129); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4131 = 8'h61 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4130); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4132 = 8'h62 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4131); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4133 = 8'h63 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4132); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4134 = 8'h64 == _T_27[7:0] ? $signed(regsA_50_re) : $signed(_GEN_4133); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4135 = 8'h65 == _T_27[7:0] ? $signed(regsA_51_re) : $signed(_GEN_4134); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4136 = 8'h66 == _T_27[7:0] ? $signed(regsA_52_re) : $signed(_GEN_4135); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4137 = 8'h67 == _T_27[7:0] ? $signed(regsA_53_re) : $signed(_GEN_4136); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4138 = 8'h68 == _T_27[7:0] ? $signed(regsA_54_re) : $signed(_GEN_4137); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4139 = 8'h69 == _T_27[7:0] ? $signed(regsA_55_re) : $signed(_GEN_4138); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4140 = 8'h6a == _T_27[7:0] ? $signed(regsA_56_re) : $signed(_GEN_4139); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4141 = 8'h6b == _T_27[7:0] ? $signed(regsA_57_re) : $signed(_GEN_4140); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4142 = 8'h6c == _T_27[7:0] ? $signed(regsA_58_re) : $signed(_GEN_4141); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4143 = 8'h6d == _T_27[7:0] ? $signed(regsA_59_re) : $signed(_GEN_4142); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4144 = 8'h6e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4143); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4145 = 8'h6f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4144); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4146 = 8'h70 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4145); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4147 = 8'h71 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4146); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4148 = 8'h72 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4147); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4149 = 8'h73 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4148); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4150 = 8'h74 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4149); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4151 = 8'h75 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4150); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4152 = 8'h76 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4151); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4153 = 8'h77 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4152); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4154 = 8'h78 == _T_27[7:0] ? $signed(regsA_60_re) : $signed(_GEN_4153); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4155 = 8'h79 == _T_27[7:0] ? $signed(regsA_61_re) : $signed(_GEN_4154); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4156 = 8'h7a == _T_27[7:0] ? $signed(regsA_62_re) : $signed(_GEN_4155); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4157 = 8'h7b == _T_27[7:0] ? $signed(regsA_63_re) : $signed(_GEN_4156); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4158 = 8'h7c == _T_27[7:0] ? $signed(regsA_64_re) : $signed(_GEN_4157); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4159 = 8'h7d == _T_27[7:0] ? $signed(regsA_65_re) : $signed(_GEN_4158); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4160 = 8'h7e == _T_27[7:0] ? $signed(regsA_66_re) : $signed(_GEN_4159); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4161 = 8'h7f == _T_27[7:0] ? $signed(regsA_67_re) : $signed(_GEN_4160); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4162 = 8'h80 == _T_27[7:0] ? $signed(regsA_68_re) : $signed(_GEN_4161); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4163 = 8'h81 == _T_27[7:0] ? $signed(regsA_69_re) : $signed(_GEN_4162); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4164 = 8'h82 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4163); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4165 = 8'h83 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4164); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4166 = 8'h84 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4165); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4167 = 8'h85 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4166); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4168 = 8'h86 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4167); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4169 = 8'h87 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4168); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4170 = 8'h88 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4169); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4171 = 8'h89 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4170); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4172 = 8'h8a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4171); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4173 = 8'h8b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4172); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4174 = 8'h8c == _T_27[7:0] ? $signed(regsA_70_re) : $signed(_GEN_4173); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4175 = 8'h8d == _T_27[7:0] ? $signed(regsA_71_re) : $signed(_GEN_4174); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4176 = 8'h8e == _T_27[7:0] ? $signed(regsA_72_re) : $signed(_GEN_4175); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4177 = 8'h8f == _T_27[7:0] ? $signed(regsA_73_re) : $signed(_GEN_4176); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4178 = 8'h90 == _T_27[7:0] ? $signed(regsA_74_re) : $signed(_GEN_4177); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4179 = 8'h91 == _T_27[7:0] ? $signed(regsA_75_re) : $signed(_GEN_4178); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4180 = 8'h92 == _T_27[7:0] ? $signed(regsA_76_re) : $signed(_GEN_4179); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4181 = 8'h93 == _T_27[7:0] ? $signed(regsA_77_re) : $signed(_GEN_4180); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4182 = 8'h94 == _T_27[7:0] ? $signed(regsA_78_re) : $signed(_GEN_4181); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4183 = 8'h95 == _T_27[7:0] ? $signed(regsA_79_re) : $signed(_GEN_4182); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4184 = 8'h96 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4183); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4185 = 8'h97 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4184); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4186 = 8'h98 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4185); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4187 = 8'h99 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4186); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4188 = 8'h9a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4187); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4189 = 8'h9b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4188); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4190 = 8'h9c == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4189); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4191 = 8'h9d == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4190); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4192 = 8'h9e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4191); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4193 = 8'h9f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4192); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4194 = 8'ha0 == _T_27[7:0] ? $signed(regsA_80_re) : $signed(_GEN_4193); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4195 = 8'ha1 == _T_27[7:0] ? $signed(regsA_81_re) : $signed(_GEN_4194); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4196 = 8'ha2 == _T_27[7:0] ? $signed(regsA_82_re) : $signed(_GEN_4195); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4197 = 8'ha3 == _T_27[7:0] ? $signed(regsA_83_re) : $signed(_GEN_4196); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4198 = 8'ha4 == _T_27[7:0] ? $signed(regsA_84_re) : $signed(_GEN_4197); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4199 = 8'ha5 == _T_27[7:0] ? $signed(regsA_85_re) : $signed(_GEN_4198); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4200 = 8'ha6 == _T_27[7:0] ? $signed(regsA_86_re) : $signed(_GEN_4199); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4201 = 8'ha7 == _T_27[7:0] ? $signed(regsA_87_re) : $signed(_GEN_4200); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4202 = 8'ha8 == _T_27[7:0] ? $signed(regsA_88_re) : $signed(_GEN_4201); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4203 = 8'ha9 == _T_27[7:0] ? $signed(regsA_89_re) : $signed(_GEN_4202); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4204 = 8'haa == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4203); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4205 = 8'hab == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4204); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4206 = 8'hac == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4205); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4207 = 8'had == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4206); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4208 = 8'hae == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4207); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4209 = 8'haf == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4208); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4210 = 8'hb0 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4209); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4211 = 8'hb1 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4210); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4212 = 8'hb2 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4211); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4213 = 8'hb3 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_4212); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4214 = 8'hb4 == _T_27[7:0] ? $signed(regsA_90_re) : $signed(_GEN_4213); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4215 = 8'hb5 == _T_27[7:0] ? $signed(regsA_91_re) : $signed(_GEN_4214); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4216 = 8'hb6 == _T_27[7:0] ? $signed(regsA_92_re) : $signed(_GEN_4215); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4217 = 8'hb7 == _T_27[7:0] ? $signed(regsA_93_re) : $signed(_GEN_4216); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4218 = 8'hb8 == _T_27[7:0] ? $signed(regsA_94_re) : $signed(_GEN_4217); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4219 = 8'hb9 == _T_27[7:0] ? $signed(regsA_95_re) : $signed(_GEN_4218); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4220 = 8'hba == _T_27[7:0] ? $signed(regsA_96_re) : $signed(_GEN_4219); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4221 = 8'hbb == _T_27[7:0] ? $signed(regsA_97_re) : $signed(_GEN_4220); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4222 = 8'hbc == _T_27[7:0] ? $signed(regsA_98_re) : $signed(_GEN_4221); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4223 = 8'hbd == _T_27[7:0] ? $signed(regsA_99_re) : $signed(_GEN_4222); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [8:0] _T_29 = 4'h9 * 5'h13; // @[Matrix_Mul_V1.scala 148:44]
  wire [8:0] _T_31 = _T_29 + _GEN_9203; // @[Matrix_Mul_V1.scala 148:60]
  wire [31:0] _GEN_4225 = 8'h1 == _T_31[7:0] ? $signed(regsA_1_im) : $signed(regsA_0_im); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4226 = 8'h2 == _T_31[7:0] ? $signed(regsA_2_im) : $signed(_GEN_4225); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4227 = 8'h3 == _T_31[7:0] ? $signed(regsA_3_im) : $signed(_GEN_4226); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4228 = 8'h4 == _T_31[7:0] ? $signed(regsA_4_im) : $signed(_GEN_4227); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4229 = 8'h5 == _T_31[7:0] ? $signed(regsA_5_im) : $signed(_GEN_4228); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4230 = 8'h6 == _T_31[7:0] ? $signed(regsA_6_im) : $signed(_GEN_4229); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4231 = 8'h7 == _T_31[7:0] ? $signed(regsA_7_im) : $signed(_GEN_4230); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4232 = 8'h8 == _T_31[7:0] ? $signed(regsA_8_im) : $signed(_GEN_4231); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4233 = 8'h9 == _T_31[7:0] ? $signed(regsA_9_im) : $signed(_GEN_4232); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4234 = 8'ha == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4233); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4235 = 8'hb == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4234); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4236 = 8'hc == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4235); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4237 = 8'hd == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4236); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4238 = 8'he == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4237); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4239 = 8'hf == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4238); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4240 = 8'h10 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4239); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4241 = 8'h11 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4240); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4242 = 8'h12 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4241); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4243 = 8'h13 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4242); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4244 = 8'h14 == _T_31[7:0] ? $signed(regsA_10_im) : $signed(_GEN_4243); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4245 = 8'h15 == _T_31[7:0] ? $signed(regsA_11_im) : $signed(_GEN_4244); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4246 = 8'h16 == _T_31[7:0] ? $signed(regsA_12_im) : $signed(_GEN_4245); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4247 = 8'h17 == _T_31[7:0] ? $signed(regsA_13_im) : $signed(_GEN_4246); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4248 = 8'h18 == _T_31[7:0] ? $signed(regsA_14_im) : $signed(_GEN_4247); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4249 = 8'h19 == _T_31[7:0] ? $signed(regsA_15_im) : $signed(_GEN_4248); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4250 = 8'h1a == _T_31[7:0] ? $signed(regsA_16_im) : $signed(_GEN_4249); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4251 = 8'h1b == _T_31[7:0] ? $signed(regsA_17_im) : $signed(_GEN_4250); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4252 = 8'h1c == _T_31[7:0] ? $signed(regsA_18_im) : $signed(_GEN_4251); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4253 = 8'h1d == _T_31[7:0] ? $signed(regsA_19_im) : $signed(_GEN_4252); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4254 = 8'h1e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4253); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4255 = 8'h1f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4254); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4256 = 8'h20 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4255); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4257 = 8'h21 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4256); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4258 = 8'h22 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4257); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4259 = 8'h23 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4258); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4260 = 8'h24 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4259); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4261 = 8'h25 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4260); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4262 = 8'h26 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4261); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4263 = 8'h27 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4262); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4264 = 8'h28 == _T_31[7:0] ? $signed(regsA_20_im) : $signed(_GEN_4263); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4265 = 8'h29 == _T_31[7:0] ? $signed(regsA_21_im) : $signed(_GEN_4264); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4266 = 8'h2a == _T_31[7:0] ? $signed(regsA_22_im) : $signed(_GEN_4265); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4267 = 8'h2b == _T_31[7:0] ? $signed(regsA_23_im) : $signed(_GEN_4266); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4268 = 8'h2c == _T_31[7:0] ? $signed(regsA_24_im) : $signed(_GEN_4267); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4269 = 8'h2d == _T_31[7:0] ? $signed(regsA_25_im) : $signed(_GEN_4268); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4270 = 8'h2e == _T_31[7:0] ? $signed(regsA_26_im) : $signed(_GEN_4269); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4271 = 8'h2f == _T_31[7:0] ? $signed(regsA_27_im) : $signed(_GEN_4270); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4272 = 8'h30 == _T_31[7:0] ? $signed(regsA_28_im) : $signed(_GEN_4271); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4273 = 8'h31 == _T_31[7:0] ? $signed(regsA_29_im) : $signed(_GEN_4272); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4274 = 8'h32 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4273); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4275 = 8'h33 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4274); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4276 = 8'h34 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4275); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4277 = 8'h35 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4276); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4278 = 8'h36 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4277); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4279 = 8'h37 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4278); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4280 = 8'h38 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4279); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4281 = 8'h39 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4280); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4282 = 8'h3a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4281); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4283 = 8'h3b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4282); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4284 = 8'h3c == _T_31[7:0] ? $signed(regsA_30_im) : $signed(_GEN_4283); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4285 = 8'h3d == _T_31[7:0] ? $signed(regsA_31_im) : $signed(_GEN_4284); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4286 = 8'h3e == _T_31[7:0] ? $signed(regsA_32_im) : $signed(_GEN_4285); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4287 = 8'h3f == _T_31[7:0] ? $signed(regsA_33_im) : $signed(_GEN_4286); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4288 = 8'h40 == _T_31[7:0] ? $signed(regsA_34_im) : $signed(_GEN_4287); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4289 = 8'h41 == _T_31[7:0] ? $signed(regsA_35_im) : $signed(_GEN_4288); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4290 = 8'h42 == _T_31[7:0] ? $signed(regsA_36_im) : $signed(_GEN_4289); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4291 = 8'h43 == _T_31[7:0] ? $signed(regsA_37_im) : $signed(_GEN_4290); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4292 = 8'h44 == _T_31[7:0] ? $signed(regsA_38_im) : $signed(_GEN_4291); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4293 = 8'h45 == _T_31[7:0] ? $signed(regsA_39_im) : $signed(_GEN_4292); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4294 = 8'h46 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4293); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4295 = 8'h47 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4294); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4296 = 8'h48 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4295); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4297 = 8'h49 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4296); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4298 = 8'h4a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4297); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4299 = 8'h4b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4298); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4300 = 8'h4c == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4299); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4301 = 8'h4d == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4300); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4302 = 8'h4e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4301); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4303 = 8'h4f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4302); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4304 = 8'h50 == _T_31[7:0] ? $signed(regsA_40_im) : $signed(_GEN_4303); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4305 = 8'h51 == _T_31[7:0] ? $signed(regsA_41_im) : $signed(_GEN_4304); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4306 = 8'h52 == _T_31[7:0] ? $signed(regsA_42_im) : $signed(_GEN_4305); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4307 = 8'h53 == _T_31[7:0] ? $signed(regsA_43_im) : $signed(_GEN_4306); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4308 = 8'h54 == _T_31[7:0] ? $signed(regsA_44_im) : $signed(_GEN_4307); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4309 = 8'h55 == _T_31[7:0] ? $signed(regsA_45_im) : $signed(_GEN_4308); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4310 = 8'h56 == _T_31[7:0] ? $signed(regsA_46_im) : $signed(_GEN_4309); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4311 = 8'h57 == _T_31[7:0] ? $signed(regsA_47_im) : $signed(_GEN_4310); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4312 = 8'h58 == _T_31[7:0] ? $signed(regsA_48_im) : $signed(_GEN_4311); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4313 = 8'h59 == _T_31[7:0] ? $signed(regsA_49_im) : $signed(_GEN_4312); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4314 = 8'h5a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4313); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4315 = 8'h5b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4314); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4316 = 8'h5c == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4315); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4317 = 8'h5d == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4316); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4318 = 8'h5e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4317); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4319 = 8'h5f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4318); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4320 = 8'h60 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4319); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4321 = 8'h61 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4320); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4322 = 8'h62 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4321); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4323 = 8'h63 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4322); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4324 = 8'h64 == _T_31[7:0] ? $signed(regsA_50_im) : $signed(_GEN_4323); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4325 = 8'h65 == _T_31[7:0] ? $signed(regsA_51_im) : $signed(_GEN_4324); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4326 = 8'h66 == _T_31[7:0] ? $signed(regsA_52_im) : $signed(_GEN_4325); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4327 = 8'h67 == _T_31[7:0] ? $signed(regsA_53_im) : $signed(_GEN_4326); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4328 = 8'h68 == _T_31[7:0] ? $signed(regsA_54_im) : $signed(_GEN_4327); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4329 = 8'h69 == _T_31[7:0] ? $signed(regsA_55_im) : $signed(_GEN_4328); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4330 = 8'h6a == _T_31[7:0] ? $signed(regsA_56_im) : $signed(_GEN_4329); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4331 = 8'h6b == _T_31[7:0] ? $signed(regsA_57_im) : $signed(_GEN_4330); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4332 = 8'h6c == _T_31[7:0] ? $signed(regsA_58_im) : $signed(_GEN_4331); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4333 = 8'h6d == _T_31[7:0] ? $signed(regsA_59_im) : $signed(_GEN_4332); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4334 = 8'h6e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4333); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4335 = 8'h6f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4334); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4336 = 8'h70 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4335); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4337 = 8'h71 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4336); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4338 = 8'h72 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4337); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4339 = 8'h73 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4338); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4340 = 8'h74 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4339); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4341 = 8'h75 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4340); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4342 = 8'h76 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4341); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4343 = 8'h77 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4342); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4344 = 8'h78 == _T_31[7:0] ? $signed(regsA_60_im) : $signed(_GEN_4343); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4345 = 8'h79 == _T_31[7:0] ? $signed(regsA_61_im) : $signed(_GEN_4344); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4346 = 8'h7a == _T_31[7:0] ? $signed(regsA_62_im) : $signed(_GEN_4345); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4347 = 8'h7b == _T_31[7:0] ? $signed(regsA_63_im) : $signed(_GEN_4346); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4348 = 8'h7c == _T_31[7:0] ? $signed(regsA_64_im) : $signed(_GEN_4347); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4349 = 8'h7d == _T_31[7:0] ? $signed(regsA_65_im) : $signed(_GEN_4348); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4350 = 8'h7e == _T_31[7:0] ? $signed(regsA_66_im) : $signed(_GEN_4349); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4351 = 8'h7f == _T_31[7:0] ? $signed(regsA_67_im) : $signed(_GEN_4350); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4352 = 8'h80 == _T_31[7:0] ? $signed(regsA_68_im) : $signed(_GEN_4351); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4353 = 8'h81 == _T_31[7:0] ? $signed(regsA_69_im) : $signed(_GEN_4352); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4354 = 8'h82 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4353); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4355 = 8'h83 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4354); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4356 = 8'h84 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4355); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4357 = 8'h85 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4356); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4358 = 8'h86 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4357); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4359 = 8'h87 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4358); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4360 = 8'h88 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4359); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4361 = 8'h89 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4360); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4362 = 8'h8a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4361); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4363 = 8'h8b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4362); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4364 = 8'h8c == _T_31[7:0] ? $signed(regsA_70_im) : $signed(_GEN_4363); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4365 = 8'h8d == _T_31[7:0] ? $signed(regsA_71_im) : $signed(_GEN_4364); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4366 = 8'h8e == _T_31[7:0] ? $signed(regsA_72_im) : $signed(_GEN_4365); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4367 = 8'h8f == _T_31[7:0] ? $signed(regsA_73_im) : $signed(_GEN_4366); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4368 = 8'h90 == _T_31[7:0] ? $signed(regsA_74_im) : $signed(_GEN_4367); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4369 = 8'h91 == _T_31[7:0] ? $signed(regsA_75_im) : $signed(_GEN_4368); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4370 = 8'h92 == _T_31[7:0] ? $signed(regsA_76_im) : $signed(_GEN_4369); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4371 = 8'h93 == _T_31[7:0] ? $signed(regsA_77_im) : $signed(_GEN_4370); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4372 = 8'h94 == _T_31[7:0] ? $signed(regsA_78_im) : $signed(_GEN_4371); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4373 = 8'h95 == _T_31[7:0] ? $signed(regsA_79_im) : $signed(_GEN_4372); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4374 = 8'h96 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4373); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4375 = 8'h97 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4374); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4376 = 8'h98 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4375); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4377 = 8'h99 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4376); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4378 = 8'h9a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4377); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4379 = 8'h9b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4378); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4380 = 8'h9c == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4379); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4381 = 8'h9d == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4380); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4382 = 8'h9e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4381); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4383 = 8'h9f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4382); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4384 = 8'ha0 == _T_31[7:0] ? $signed(regsA_80_im) : $signed(_GEN_4383); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4385 = 8'ha1 == _T_31[7:0] ? $signed(regsA_81_im) : $signed(_GEN_4384); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4386 = 8'ha2 == _T_31[7:0] ? $signed(regsA_82_im) : $signed(_GEN_4385); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4387 = 8'ha3 == _T_31[7:0] ? $signed(regsA_83_im) : $signed(_GEN_4386); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4388 = 8'ha4 == _T_31[7:0] ? $signed(regsA_84_im) : $signed(_GEN_4387); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4389 = 8'ha5 == _T_31[7:0] ? $signed(regsA_85_im) : $signed(_GEN_4388); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4390 = 8'ha6 == _T_31[7:0] ? $signed(regsA_86_im) : $signed(_GEN_4389); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4391 = 8'ha7 == _T_31[7:0] ? $signed(regsA_87_im) : $signed(_GEN_4390); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4392 = 8'ha8 == _T_31[7:0] ? $signed(regsA_88_im) : $signed(_GEN_4391); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4393 = 8'ha9 == _T_31[7:0] ? $signed(regsA_89_im) : $signed(_GEN_4392); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4394 = 8'haa == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4393); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4395 = 8'hab == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4394); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4396 = 8'hac == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4395); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4397 = 8'had == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4396); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4398 = 8'hae == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4397); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4399 = 8'haf == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4398); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4400 = 8'hb0 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4399); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4401 = 8'hb1 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4400); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4402 = 8'hb2 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4401); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4403 = 8'hb3 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4402); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4404 = 8'hb4 == _T_31[7:0] ? $signed(regsA_90_im) : $signed(_GEN_4403); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4405 = 8'hb5 == _T_31[7:0] ? $signed(regsA_91_im) : $signed(_GEN_4404); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4406 = 8'hb6 == _T_31[7:0] ? $signed(regsA_92_im) : $signed(_GEN_4405); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4407 = 8'hb7 == _T_31[7:0] ? $signed(regsA_93_im) : $signed(_GEN_4406); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4408 = 8'hb8 == _T_31[7:0] ? $signed(regsA_94_im) : $signed(_GEN_4407); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4409 = 8'hb9 == _T_31[7:0] ? $signed(regsA_95_im) : $signed(_GEN_4408); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4410 = 8'hba == _T_31[7:0] ? $signed(regsA_96_im) : $signed(_GEN_4409); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4411 = 8'hbb == _T_31[7:0] ? $signed(regsA_97_im) : $signed(_GEN_4410); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4412 = 8'hbc == _T_31[7:0] ? $signed(regsA_98_im) : $signed(_GEN_4411); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4413 = 8'hbd == _T_31[7:0] ? $signed(regsA_99_im) : $signed(_GEN_4412); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4415 = 8'h1 == _T_31[7:0] ? $signed(regsA_1_re) : $signed(regsA_0_re); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4416 = 8'h2 == _T_31[7:0] ? $signed(regsA_2_re) : $signed(_GEN_4415); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4417 = 8'h3 == _T_31[7:0] ? $signed(regsA_3_re) : $signed(_GEN_4416); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4418 = 8'h4 == _T_31[7:0] ? $signed(regsA_4_re) : $signed(_GEN_4417); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4419 = 8'h5 == _T_31[7:0] ? $signed(regsA_5_re) : $signed(_GEN_4418); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4420 = 8'h6 == _T_31[7:0] ? $signed(regsA_6_re) : $signed(_GEN_4419); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4421 = 8'h7 == _T_31[7:0] ? $signed(regsA_7_re) : $signed(_GEN_4420); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4422 = 8'h8 == _T_31[7:0] ? $signed(regsA_8_re) : $signed(_GEN_4421); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4423 = 8'h9 == _T_31[7:0] ? $signed(regsA_9_re) : $signed(_GEN_4422); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4424 = 8'ha == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4423); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4425 = 8'hb == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4424); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4426 = 8'hc == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4425); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4427 = 8'hd == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4426); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4428 = 8'he == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4427); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4429 = 8'hf == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4428); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4430 = 8'h10 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4429); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4431 = 8'h11 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4430); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4432 = 8'h12 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4431); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4433 = 8'h13 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4432); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4434 = 8'h14 == _T_31[7:0] ? $signed(regsA_10_re) : $signed(_GEN_4433); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4435 = 8'h15 == _T_31[7:0] ? $signed(regsA_11_re) : $signed(_GEN_4434); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4436 = 8'h16 == _T_31[7:0] ? $signed(regsA_12_re) : $signed(_GEN_4435); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4437 = 8'h17 == _T_31[7:0] ? $signed(regsA_13_re) : $signed(_GEN_4436); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4438 = 8'h18 == _T_31[7:0] ? $signed(regsA_14_re) : $signed(_GEN_4437); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4439 = 8'h19 == _T_31[7:0] ? $signed(regsA_15_re) : $signed(_GEN_4438); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4440 = 8'h1a == _T_31[7:0] ? $signed(regsA_16_re) : $signed(_GEN_4439); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4441 = 8'h1b == _T_31[7:0] ? $signed(regsA_17_re) : $signed(_GEN_4440); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4442 = 8'h1c == _T_31[7:0] ? $signed(regsA_18_re) : $signed(_GEN_4441); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4443 = 8'h1d == _T_31[7:0] ? $signed(regsA_19_re) : $signed(_GEN_4442); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4444 = 8'h1e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4443); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4445 = 8'h1f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4444); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4446 = 8'h20 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4445); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4447 = 8'h21 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4446); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4448 = 8'h22 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4447); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4449 = 8'h23 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4448); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4450 = 8'h24 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4449); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4451 = 8'h25 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4450); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4452 = 8'h26 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4451); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4453 = 8'h27 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4452); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4454 = 8'h28 == _T_31[7:0] ? $signed(regsA_20_re) : $signed(_GEN_4453); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4455 = 8'h29 == _T_31[7:0] ? $signed(regsA_21_re) : $signed(_GEN_4454); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4456 = 8'h2a == _T_31[7:0] ? $signed(regsA_22_re) : $signed(_GEN_4455); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4457 = 8'h2b == _T_31[7:0] ? $signed(regsA_23_re) : $signed(_GEN_4456); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4458 = 8'h2c == _T_31[7:0] ? $signed(regsA_24_re) : $signed(_GEN_4457); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4459 = 8'h2d == _T_31[7:0] ? $signed(regsA_25_re) : $signed(_GEN_4458); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4460 = 8'h2e == _T_31[7:0] ? $signed(regsA_26_re) : $signed(_GEN_4459); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4461 = 8'h2f == _T_31[7:0] ? $signed(regsA_27_re) : $signed(_GEN_4460); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4462 = 8'h30 == _T_31[7:0] ? $signed(regsA_28_re) : $signed(_GEN_4461); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4463 = 8'h31 == _T_31[7:0] ? $signed(regsA_29_re) : $signed(_GEN_4462); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4464 = 8'h32 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4463); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4465 = 8'h33 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4464); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4466 = 8'h34 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4465); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4467 = 8'h35 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4466); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4468 = 8'h36 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4467); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4469 = 8'h37 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4468); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4470 = 8'h38 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4469); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4471 = 8'h39 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4470); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4472 = 8'h3a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4471); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4473 = 8'h3b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4472); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4474 = 8'h3c == _T_31[7:0] ? $signed(regsA_30_re) : $signed(_GEN_4473); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4475 = 8'h3d == _T_31[7:0] ? $signed(regsA_31_re) : $signed(_GEN_4474); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4476 = 8'h3e == _T_31[7:0] ? $signed(regsA_32_re) : $signed(_GEN_4475); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4477 = 8'h3f == _T_31[7:0] ? $signed(regsA_33_re) : $signed(_GEN_4476); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4478 = 8'h40 == _T_31[7:0] ? $signed(regsA_34_re) : $signed(_GEN_4477); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4479 = 8'h41 == _T_31[7:0] ? $signed(regsA_35_re) : $signed(_GEN_4478); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4480 = 8'h42 == _T_31[7:0] ? $signed(regsA_36_re) : $signed(_GEN_4479); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4481 = 8'h43 == _T_31[7:0] ? $signed(regsA_37_re) : $signed(_GEN_4480); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4482 = 8'h44 == _T_31[7:0] ? $signed(regsA_38_re) : $signed(_GEN_4481); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4483 = 8'h45 == _T_31[7:0] ? $signed(regsA_39_re) : $signed(_GEN_4482); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4484 = 8'h46 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4483); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4485 = 8'h47 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4484); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4486 = 8'h48 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4485); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4487 = 8'h49 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4486); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4488 = 8'h4a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4487); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4489 = 8'h4b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4488); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4490 = 8'h4c == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4489); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4491 = 8'h4d == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4490); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4492 = 8'h4e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4491); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4493 = 8'h4f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4492); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4494 = 8'h50 == _T_31[7:0] ? $signed(regsA_40_re) : $signed(_GEN_4493); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4495 = 8'h51 == _T_31[7:0] ? $signed(regsA_41_re) : $signed(_GEN_4494); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4496 = 8'h52 == _T_31[7:0] ? $signed(regsA_42_re) : $signed(_GEN_4495); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4497 = 8'h53 == _T_31[7:0] ? $signed(regsA_43_re) : $signed(_GEN_4496); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4498 = 8'h54 == _T_31[7:0] ? $signed(regsA_44_re) : $signed(_GEN_4497); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4499 = 8'h55 == _T_31[7:0] ? $signed(regsA_45_re) : $signed(_GEN_4498); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4500 = 8'h56 == _T_31[7:0] ? $signed(regsA_46_re) : $signed(_GEN_4499); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4501 = 8'h57 == _T_31[7:0] ? $signed(regsA_47_re) : $signed(_GEN_4500); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4502 = 8'h58 == _T_31[7:0] ? $signed(regsA_48_re) : $signed(_GEN_4501); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4503 = 8'h59 == _T_31[7:0] ? $signed(regsA_49_re) : $signed(_GEN_4502); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4504 = 8'h5a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4503); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4505 = 8'h5b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4504); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4506 = 8'h5c == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4505); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4507 = 8'h5d == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4506); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4508 = 8'h5e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4507); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4509 = 8'h5f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4508); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4510 = 8'h60 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4509); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4511 = 8'h61 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4510); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4512 = 8'h62 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4511); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4513 = 8'h63 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4512); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4514 = 8'h64 == _T_31[7:0] ? $signed(regsA_50_re) : $signed(_GEN_4513); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4515 = 8'h65 == _T_31[7:0] ? $signed(regsA_51_re) : $signed(_GEN_4514); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4516 = 8'h66 == _T_31[7:0] ? $signed(regsA_52_re) : $signed(_GEN_4515); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4517 = 8'h67 == _T_31[7:0] ? $signed(regsA_53_re) : $signed(_GEN_4516); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4518 = 8'h68 == _T_31[7:0] ? $signed(regsA_54_re) : $signed(_GEN_4517); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4519 = 8'h69 == _T_31[7:0] ? $signed(regsA_55_re) : $signed(_GEN_4518); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4520 = 8'h6a == _T_31[7:0] ? $signed(regsA_56_re) : $signed(_GEN_4519); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4521 = 8'h6b == _T_31[7:0] ? $signed(regsA_57_re) : $signed(_GEN_4520); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4522 = 8'h6c == _T_31[7:0] ? $signed(regsA_58_re) : $signed(_GEN_4521); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4523 = 8'h6d == _T_31[7:0] ? $signed(regsA_59_re) : $signed(_GEN_4522); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4524 = 8'h6e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4523); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4525 = 8'h6f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4524); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4526 = 8'h70 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4525); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4527 = 8'h71 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4526); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4528 = 8'h72 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4527); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4529 = 8'h73 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4528); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4530 = 8'h74 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4529); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4531 = 8'h75 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4530); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4532 = 8'h76 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4531); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4533 = 8'h77 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4532); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4534 = 8'h78 == _T_31[7:0] ? $signed(regsA_60_re) : $signed(_GEN_4533); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4535 = 8'h79 == _T_31[7:0] ? $signed(regsA_61_re) : $signed(_GEN_4534); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4536 = 8'h7a == _T_31[7:0] ? $signed(regsA_62_re) : $signed(_GEN_4535); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4537 = 8'h7b == _T_31[7:0] ? $signed(regsA_63_re) : $signed(_GEN_4536); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4538 = 8'h7c == _T_31[7:0] ? $signed(regsA_64_re) : $signed(_GEN_4537); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4539 = 8'h7d == _T_31[7:0] ? $signed(regsA_65_re) : $signed(_GEN_4538); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4540 = 8'h7e == _T_31[7:0] ? $signed(regsA_66_re) : $signed(_GEN_4539); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4541 = 8'h7f == _T_31[7:0] ? $signed(regsA_67_re) : $signed(_GEN_4540); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4542 = 8'h80 == _T_31[7:0] ? $signed(regsA_68_re) : $signed(_GEN_4541); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4543 = 8'h81 == _T_31[7:0] ? $signed(regsA_69_re) : $signed(_GEN_4542); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4544 = 8'h82 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4543); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4545 = 8'h83 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4544); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4546 = 8'h84 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4545); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4547 = 8'h85 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4546); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4548 = 8'h86 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4547); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4549 = 8'h87 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4548); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4550 = 8'h88 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4549); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4551 = 8'h89 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4550); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4552 = 8'h8a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4551); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4553 = 8'h8b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4552); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4554 = 8'h8c == _T_31[7:0] ? $signed(regsA_70_re) : $signed(_GEN_4553); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4555 = 8'h8d == _T_31[7:0] ? $signed(regsA_71_re) : $signed(_GEN_4554); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4556 = 8'h8e == _T_31[7:0] ? $signed(regsA_72_re) : $signed(_GEN_4555); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4557 = 8'h8f == _T_31[7:0] ? $signed(regsA_73_re) : $signed(_GEN_4556); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4558 = 8'h90 == _T_31[7:0] ? $signed(regsA_74_re) : $signed(_GEN_4557); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4559 = 8'h91 == _T_31[7:0] ? $signed(regsA_75_re) : $signed(_GEN_4558); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4560 = 8'h92 == _T_31[7:0] ? $signed(regsA_76_re) : $signed(_GEN_4559); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4561 = 8'h93 == _T_31[7:0] ? $signed(regsA_77_re) : $signed(_GEN_4560); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4562 = 8'h94 == _T_31[7:0] ? $signed(regsA_78_re) : $signed(_GEN_4561); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4563 = 8'h95 == _T_31[7:0] ? $signed(regsA_79_re) : $signed(_GEN_4562); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4564 = 8'h96 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4563); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4565 = 8'h97 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4564); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4566 = 8'h98 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4565); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4567 = 8'h99 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4566); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4568 = 8'h9a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4567); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4569 = 8'h9b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4568); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4570 = 8'h9c == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4569); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4571 = 8'h9d == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4570); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4572 = 8'h9e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4571); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4573 = 8'h9f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4572); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4574 = 8'ha0 == _T_31[7:0] ? $signed(regsA_80_re) : $signed(_GEN_4573); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4575 = 8'ha1 == _T_31[7:0] ? $signed(regsA_81_re) : $signed(_GEN_4574); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4576 = 8'ha2 == _T_31[7:0] ? $signed(regsA_82_re) : $signed(_GEN_4575); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4577 = 8'ha3 == _T_31[7:0] ? $signed(regsA_83_re) : $signed(_GEN_4576); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4578 = 8'ha4 == _T_31[7:0] ? $signed(regsA_84_re) : $signed(_GEN_4577); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4579 = 8'ha5 == _T_31[7:0] ? $signed(regsA_85_re) : $signed(_GEN_4578); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4580 = 8'ha6 == _T_31[7:0] ? $signed(regsA_86_re) : $signed(_GEN_4579); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4581 = 8'ha7 == _T_31[7:0] ? $signed(regsA_87_re) : $signed(_GEN_4580); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4582 = 8'ha8 == _T_31[7:0] ? $signed(regsA_88_re) : $signed(_GEN_4581); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4583 = 8'ha9 == _T_31[7:0] ? $signed(regsA_89_re) : $signed(_GEN_4582); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4584 = 8'haa == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4583); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4585 = 8'hab == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4584); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4586 = 8'hac == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4585); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4587 = 8'had == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4586); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4588 = 8'hae == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4587); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4589 = 8'haf == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4588); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4590 = 8'hb0 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4589); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4591 = 8'hb1 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4590); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4592 = 8'hb2 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4591); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4593 = 8'hb3 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_4592); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4594 = 8'hb4 == _T_31[7:0] ? $signed(regsA_90_re) : $signed(_GEN_4593); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4595 = 8'hb5 == _T_31[7:0] ? $signed(regsA_91_re) : $signed(_GEN_4594); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4596 = 8'hb6 == _T_31[7:0] ? $signed(regsA_92_re) : $signed(_GEN_4595); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4597 = 8'hb7 == _T_31[7:0] ? $signed(regsA_93_re) : $signed(_GEN_4596); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4598 = 8'hb8 == _T_31[7:0] ? $signed(regsA_94_re) : $signed(_GEN_4597); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4599 = 8'hb9 == _T_31[7:0] ? $signed(regsA_95_re) : $signed(_GEN_4598); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4600 = 8'hba == _T_31[7:0] ? $signed(regsA_96_re) : $signed(_GEN_4599); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4601 = 8'hbb == _T_31[7:0] ? $signed(regsA_97_re) : $signed(_GEN_4600); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4602 = 8'hbc == _T_31[7:0] ? $signed(regsA_98_re) : $signed(_GEN_4601); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4603 = 8'hbd == _T_31[7:0] ? $signed(regsA_99_re) : $signed(_GEN_4602); // @[Matrix_Mul_V1.scala 148:{27,27}]
  wire [31:0] _GEN_4625 = 6'h1 == _T_3 ? $signed(regsB_10_im) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4626 = 6'h2 == _T_3 ? $signed(regsB_20_im) : $signed(_GEN_4625); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4627 = 6'h3 == _T_3 ? $signed(regsB_30_im) : $signed(_GEN_4626); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4628 = 6'h4 == _T_3 ? $signed(regsB_40_im) : $signed(_GEN_4627); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4629 = 6'h5 == _T_3 ? $signed(regsB_50_im) : $signed(_GEN_4628); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4630 = 6'h6 == _T_3 ? $signed(regsB_60_im) : $signed(_GEN_4629); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4631 = 6'h7 == _T_3 ? $signed(regsB_70_im) : $signed(_GEN_4630); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4632 = 6'h8 == _T_3 ? $signed(regsB_80_im) : $signed(_GEN_4631); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4633 = 6'h9 == _T_3 ? $signed(regsB_90_im) : $signed(_GEN_4632); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4634 = 6'ha == _T_3 ? $signed(32'sh0) : $signed(_GEN_4633); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4635 = 6'hb == _T_3 ? $signed(32'sh0) : $signed(_GEN_4634); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4636 = 6'hc == _T_3 ? $signed(32'sh0) : $signed(_GEN_4635); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4637 = 6'hd == _T_3 ? $signed(32'sh0) : $signed(_GEN_4636); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4638 = 6'he == _T_3 ? $signed(32'sh0) : $signed(_GEN_4637); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4639 = 6'hf == _T_3 ? $signed(32'sh0) : $signed(_GEN_4638); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4640 = 6'h10 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4639); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4641 = 6'h11 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4640); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4642 = 6'h12 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4641); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4643 = 6'h13 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4642); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4644 = 6'h14 == _T_3 ? $signed(regsB_1_im) : $signed(_GEN_4643); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4645 = 6'h15 == _T_3 ? $signed(regsB_11_im) : $signed(_GEN_4644); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4646 = 6'h16 == _T_3 ? $signed(regsB_21_im) : $signed(_GEN_4645); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4647 = 6'h17 == _T_3 ? $signed(regsB_31_im) : $signed(_GEN_4646); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4648 = 6'h18 == _T_3 ? $signed(regsB_41_im) : $signed(_GEN_4647); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4649 = 6'h19 == _T_3 ? $signed(regsB_51_im) : $signed(_GEN_4648); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4650 = 6'h1a == _T_3 ? $signed(regsB_61_im) : $signed(_GEN_4649); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4651 = 6'h1b == _T_3 ? $signed(regsB_71_im) : $signed(_GEN_4650); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4652 = 6'h1c == _T_3 ? $signed(regsB_81_im) : $signed(_GEN_4651); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4653 = 6'h1d == _T_3 ? $signed(regsB_91_im) : $signed(_GEN_4652); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4654 = 6'h1e == _T_3 ? $signed(32'sh0) : $signed(_GEN_4653); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4655 = 6'h1f == _T_3 ? $signed(32'sh0) : $signed(_GEN_4654); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4656 = 6'h20 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4655); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4657 = 6'h21 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4656); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4658 = 6'h22 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4657); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4659 = 6'h23 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4658); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4660 = 6'h24 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4659); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4661 = 6'h25 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4660); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4662 = 6'h26 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4661); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4663 = 6'h27 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4662); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4664 = 6'h28 == _T_3 ? $signed(regsB_2_im) : $signed(_GEN_4663); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4665 = 6'h29 == _T_3 ? $signed(regsB_12_im) : $signed(_GEN_4664); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4666 = 6'h2a == _T_3 ? $signed(regsB_22_im) : $signed(_GEN_4665); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4667 = 6'h2b == _T_3 ? $signed(regsB_32_im) : $signed(_GEN_4666); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4668 = 6'h2c == _T_3 ? $signed(regsB_42_im) : $signed(_GEN_4667); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4669 = 6'h2d == _T_3 ? $signed(regsB_52_im) : $signed(_GEN_4668); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4670 = 6'h2e == _T_3 ? $signed(regsB_62_im) : $signed(_GEN_4669); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4671 = 6'h2f == _T_3 ? $signed(regsB_72_im) : $signed(_GEN_4670); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4672 = 6'h30 == _T_3 ? $signed(regsB_82_im) : $signed(_GEN_4671); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4673 = 6'h31 == _T_3 ? $signed(regsB_92_im) : $signed(_GEN_4672); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4674 = 6'h32 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4673); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4675 = 6'h33 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4674); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4676 = 6'h34 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4675); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4677 = 6'h35 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4676); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4678 = 6'h36 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4677); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4679 = 6'h37 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4678); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4680 = 6'h38 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4679); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4681 = 6'h39 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4680); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4682 = 6'h3a == _T_3 ? $signed(32'sh0) : $signed(_GEN_4681); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4683 = 6'h3b == _T_3 ? $signed(32'sh0) : $signed(_GEN_4682); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4684 = 6'h3c == _T_3 ? $signed(regsB_3_im) : $signed(_GEN_4683); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4685 = 6'h3d == _T_3 ? $signed(regsB_13_im) : $signed(_GEN_4684); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4686 = 6'h3e == _T_3 ? $signed(regsB_23_im) : $signed(_GEN_4685); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4687 = 6'h3f == _T_3 ? $signed(regsB_33_im) : $signed(_GEN_4686); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4688 = 7'h40 == _GEN_8445 ? $signed(regsB_43_im) : $signed(_GEN_4687); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4689 = 7'h41 == _GEN_8445 ? $signed(regsB_53_im) : $signed(_GEN_4688); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4690 = 7'h42 == _GEN_8445 ? $signed(regsB_63_im) : $signed(_GEN_4689); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4691 = 7'h43 == _GEN_8445 ? $signed(regsB_73_im) : $signed(_GEN_4690); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4692 = 7'h44 == _GEN_8445 ? $signed(regsB_83_im) : $signed(_GEN_4691); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4693 = 7'h45 == _GEN_8445 ? $signed(regsB_93_im) : $signed(_GEN_4692); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4694 = 7'h46 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4693); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4695 = 7'h47 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4694); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4696 = 7'h48 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4695); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4697 = 7'h49 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4696); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4698 = 7'h4a == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4697); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4699 = 7'h4b == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4698); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4700 = 7'h4c == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4699); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4701 = 7'h4d == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4700); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4702 = 7'h4e == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4701); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4703 = 7'h4f == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4702); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4704 = 7'h50 == _GEN_8445 ? $signed(regsB_4_im) : $signed(_GEN_4703); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4705 = 7'h51 == _GEN_8445 ? $signed(regsB_14_im) : $signed(_GEN_4704); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4706 = 7'h52 == _GEN_8445 ? $signed(regsB_24_im) : $signed(_GEN_4705); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4707 = 7'h53 == _GEN_8445 ? $signed(regsB_34_im) : $signed(_GEN_4706); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4708 = 7'h54 == _GEN_8445 ? $signed(regsB_44_im) : $signed(_GEN_4707); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4709 = 7'h55 == _GEN_8445 ? $signed(regsB_54_im) : $signed(_GEN_4708); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4710 = 7'h56 == _GEN_8445 ? $signed(regsB_64_im) : $signed(_GEN_4709); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4711 = 7'h57 == _GEN_8445 ? $signed(regsB_74_im) : $signed(_GEN_4710); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4712 = 7'h58 == _GEN_8445 ? $signed(regsB_84_im) : $signed(_GEN_4711); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4713 = 7'h59 == _GEN_8445 ? $signed(regsB_94_im) : $signed(_GEN_4712); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4714 = 7'h5a == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4713); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4715 = 7'h5b == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4714); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4716 = 7'h5c == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4715); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4717 = 7'h5d == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4716); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4718 = 7'h5e == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4717); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4719 = 7'h5f == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4718); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4720 = 7'h60 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4719); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4721 = 7'h61 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4720); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4722 = 7'h62 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4721); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4723 = 7'h63 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4722); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4724 = 7'h64 == _GEN_8445 ? $signed(regsB_5_im) : $signed(_GEN_4723); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4725 = 7'h65 == _GEN_8445 ? $signed(regsB_15_im) : $signed(_GEN_4724); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4726 = 7'h66 == _GEN_8445 ? $signed(regsB_25_im) : $signed(_GEN_4725); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4727 = 7'h67 == _GEN_8445 ? $signed(regsB_35_im) : $signed(_GEN_4726); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4728 = 7'h68 == _GEN_8445 ? $signed(regsB_45_im) : $signed(_GEN_4727); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4729 = 7'h69 == _GEN_8445 ? $signed(regsB_55_im) : $signed(_GEN_4728); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4730 = 7'h6a == _GEN_8445 ? $signed(regsB_65_im) : $signed(_GEN_4729); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4731 = 7'h6b == _GEN_8445 ? $signed(regsB_75_im) : $signed(_GEN_4730); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4732 = 7'h6c == _GEN_8445 ? $signed(regsB_85_im) : $signed(_GEN_4731); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4733 = 7'h6d == _GEN_8445 ? $signed(regsB_95_im) : $signed(_GEN_4732); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4734 = 7'h6e == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4733); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4735 = 7'h6f == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4734); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4736 = 7'h70 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4735); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4737 = 7'h71 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4736); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4738 = 7'h72 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4737); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4739 = 7'h73 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4738); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4740 = 7'h74 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4739); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4741 = 7'h75 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4740); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4742 = 7'h76 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4741); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4743 = 7'h77 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4742); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4744 = 7'h78 == _GEN_8445 ? $signed(regsB_6_im) : $signed(_GEN_4743); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4745 = 7'h79 == _GEN_8445 ? $signed(regsB_16_im) : $signed(_GEN_4744); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4746 = 7'h7a == _GEN_8445 ? $signed(regsB_26_im) : $signed(_GEN_4745); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4747 = 7'h7b == _GEN_8445 ? $signed(regsB_36_im) : $signed(_GEN_4746); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4748 = 7'h7c == _GEN_8445 ? $signed(regsB_46_im) : $signed(_GEN_4747); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4749 = 7'h7d == _GEN_8445 ? $signed(regsB_56_im) : $signed(_GEN_4748); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4750 = 7'h7e == _GEN_8445 ? $signed(regsB_66_im) : $signed(_GEN_4749); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4751 = 7'h7f == _GEN_8445 ? $signed(regsB_76_im) : $signed(_GEN_4750); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4752 = 8'h80 == _GEN_8509 ? $signed(regsB_86_im) : $signed(_GEN_4751); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4753 = 8'h81 == _GEN_8509 ? $signed(regsB_96_im) : $signed(_GEN_4752); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4754 = 8'h82 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4753); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4755 = 8'h83 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4754); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4756 = 8'h84 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4755); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4757 = 8'h85 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4756); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4758 = 8'h86 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4757); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4759 = 8'h87 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4758); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4760 = 8'h88 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4759); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4761 = 8'h89 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4760); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4762 = 8'h8a == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4761); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4763 = 8'h8b == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4762); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4764 = 8'h8c == _GEN_8509 ? $signed(regsB_7_im) : $signed(_GEN_4763); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4765 = 8'h8d == _GEN_8509 ? $signed(regsB_17_im) : $signed(_GEN_4764); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4766 = 8'h8e == _GEN_8509 ? $signed(regsB_27_im) : $signed(_GEN_4765); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4767 = 8'h8f == _GEN_8509 ? $signed(regsB_37_im) : $signed(_GEN_4766); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4768 = 8'h90 == _GEN_8509 ? $signed(regsB_47_im) : $signed(_GEN_4767); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4769 = 8'h91 == _GEN_8509 ? $signed(regsB_57_im) : $signed(_GEN_4768); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4770 = 8'h92 == _GEN_8509 ? $signed(regsB_67_im) : $signed(_GEN_4769); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4771 = 8'h93 == _GEN_8509 ? $signed(regsB_77_im) : $signed(_GEN_4770); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4772 = 8'h94 == _GEN_8509 ? $signed(regsB_87_im) : $signed(_GEN_4771); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4773 = 8'h95 == _GEN_8509 ? $signed(regsB_97_im) : $signed(_GEN_4772); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4774 = 8'h96 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4773); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4775 = 8'h97 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4774); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4776 = 8'h98 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4775); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4777 = 8'h99 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4776); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4778 = 8'h9a == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4777); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4779 = 8'h9b == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4778); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4780 = 8'h9c == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4779); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4781 = 8'h9d == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4780); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4782 = 8'h9e == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4781); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4783 = 8'h9f == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4782); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4784 = 8'ha0 == _GEN_8509 ? $signed(regsB_8_im) : $signed(_GEN_4783); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4785 = 8'ha1 == _GEN_8509 ? $signed(regsB_18_im) : $signed(_GEN_4784); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4786 = 8'ha2 == _GEN_8509 ? $signed(regsB_28_im) : $signed(_GEN_4785); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4787 = 8'ha3 == _GEN_8509 ? $signed(regsB_38_im) : $signed(_GEN_4786); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4788 = 8'ha4 == _GEN_8509 ? $signed(regsB_48_im) : $signed(_GEN_4787); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4789 = 8'ha5 == _GEN_8509 ? $signed(regsB_58_im) : $signed(_GEN_4788); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4790 = 8'ha6 == _GEN_8509 ? $signed(regsB_68_im) : $signed(_GEN_4789); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4791 = 8'ha7 == _GEN_8509 ? $signed(regsB_78_im) : $signed(_GEN_4790); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4792 = 8'ha8 == _GEN_8509 ? $signed(regsB_88_im) : $signed(_GEN_4791); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4793 = 8'ha9 == _GEN_8509 ? $signed(regsB_98_im) : $signed(_GEN_4792); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4794 = 8'haa == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4793); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4795 = 8'hab == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4794); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4796 = 8'hac == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4795); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4797 = 8'had == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4796); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4798 = 8'hae == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4797); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4799 = 8'haf == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4798); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4800 = 8'hb0 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4799); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4801 = 8'hb1 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4800); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4802 = 8'hb2 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4801); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4803 = 8'hb3 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4802); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4804 = 8'hb4 == _GEN_8509 ? $signed(regsB_9_im) : $signed(_GEN_4803); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4805 = 8'hb5 == _GEN_8509 ? $signed(regsB_19_im) : $signed(_GEN_4804); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4806 = 8'hb6 == _GEN_8509 ? $signed(regsB_29_im) : $signed(_GEN_4805); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4807 = 8'hb7 == _GEN_8509 ? $signed(regsB_39_im) : $signed(_GEN_4806); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4808 = 8'hb8 == _GEN_8509 ? $signed(regsB_49_im) : $signed(_GEN_4807); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4809 = 8'hb9 == _GEN_8509 ? $signed(regsB_59_im) : $signed(_GEN_4808); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4810 = 8'hba == _GEN_8509 ? $signed(regsB_69_im) : $signed(_GEN_4809); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4811 = 8'hbb == _GEN_8509 ? $signed(regsB_79_im) : $signed(_GEN_4810); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4812 = 8'hbc == _GEN_8509 ? $signed(regsB_89_im) : $signed(_GEN_4811); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4813 = 8'hbd == _GEN_8509 ? $signed(regsB_99_im) : $signed(_GEN_4812); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4815 = 6'h1 == _T_3 ? $signed(regsB_10_re) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4816 = 6'h2 == _T_3 ? $signed(regsB_20_re) : $signed(_GEN_4815); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4817 = 6'h3 == _T_3 ? $signed(regsB_30_re) : $signed(_GEN_4816); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4818 = 6'h4 == _T_3 ? $signed(regsB_40_re) : $signed(_GEN_4817); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4819 = 6'h5 == _T_3 ? $signed(regsB_50_re) : $signed(_GEN_4818); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4820 = 6'h6 == _T_3 ? $signed(regsB_60_re) : $signed(_GEN_4819); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4821 = 6'h7 == _T_3 ? $signed(regsB_70_re) : $signed(_GEN_4820); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4822 = 6'h8 == _T_3 ? $signed(regsB_80_re) : $signed(_GEN_4821); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4823 = 6'h9 == _T_3 ? $signed(regsB_90_re) : $signed(_GEN_4822); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4824 = 6'ha == _T_3 ? $signed(32'sh0) : $signed(_GEN_4823); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4825 = 6'hb == _T_3 ? $signed(32'sh0) : $signed(_GEN_4824); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4826 = 6'hc == _T_3 ? $signed(32'sh0) : $signed(_GEN_4825); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4827 = 6'hd == _T_3 ? $signed(32'sh0) : $signed(_GEN_4826); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4828 = 6'he == _T_3 ? $signed(32'sh0) : $signed(_GEN_4827); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4829 = 6'hf == _T_3 ? $signed(32'sh0) : $signed(_GEN_4828); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4830 = 6'h10 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4829); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4831 = 6'h11 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4830); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4832 = 6'h12 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4831); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4833 = 6'h13 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4832); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4834 = 6'h14 == _T_3 ? $signed(regsB_1_re) : $signed(_GEN_4833); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4835 = 6'h15 == _T_3 ? $signed(regsB_11_re) : $signed(_GEN_4834); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4836 = 6'h16 == _T_3 ? $signed(regsB_21_re) : $signed(_GEN_4835); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4837 = 6'h17 == _T_3 ? $signed(regsB_31_re) : $signed(_GEN_4836); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4838 = 6'h18 == _T_3 ? $signed(regsB_41_re) : $signed(_GEN_4837); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4839 = 6'h19 == _T_3 ? $signed(regsB_51_re) : $signed(_GEN_4838); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4840 = 6'h1a == _T_3 ? $signed(regsB_61_re) : $signed(_GEN_4839); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4841 = 6'h1b == _T_3 ? $signed(regsB_71_re) : $signed(_GEN_4840); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4842 = 6'h1c == _T_3 ? $signed(regsB_81_re) : $signed(_GEN_4841); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4843 = 6'h1d == _T_3 ? $signed(regsB_91_re) : $signed(_GEN_4842); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4844 = 6'h1e == _T_3 ? $signed(32'sh0) : $signed(_GEN_4843); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4845 = 6'h1f == _T_3 ? $signed(32'sh0) : $signed(_GEN_4844); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4846 = 6'h20 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4845); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4847 = 6'h21 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4846); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4848 = 6'h22 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4847); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4849 = 6'h23 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4848); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4850 = 6'h24 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4849); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4851 = 6'h25 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4850); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4852 = 6'h26 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4851); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4853 = 6'h27 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4852); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4854 = 6'h28 == _T_3 ? $signed(regsB_2_re) : $signed(_GEN_4853); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4855 = 6'h29 == _T_3 ? $signed(regsB_12_re) : $signed(_GEN_4854); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4856 = 6'h2a == _T_3 ? $signed(regsB_22_re) : $signed(_GEN_4855); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4857 = 6'h2b == _T_3 ? $signed(regsB_32_re) : $signed(_GEN_4856); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4858 = 6'h2c == _T_3 ? $signed(regsB_42_re) : $signed(_GEN_4857); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4859 = 6'h2d == _T_3 ? $signed(regsB_52_re) : $signed(_GEN_4858); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4860 = 6'h2e == _T_3 ? $signed(regsB_62_re) : $signed(_GEN_4859); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4861 = 6'h2f == _T_3 ? $signed(regsB_72_re) : $signed(_GEN_4860); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4862 = 6'h30 == _T_3 ? $signed(regsB_82_re) : $signed(_GEN_4861); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4863 = 6'h31 == _T_3 ? $signed(regsB_92_re) : $signed(_GEN_4862); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4864 = 6'h32 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4863); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4865 = 6'h33 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4864); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4866 = 6'h34 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4865); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4867 = 6'h35 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4866); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4868 = 6'h36 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4867); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4869 = 6'h37 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4868); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4870 = 6'h38 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4869); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4871 = 6'h39 == _T_3 ? $signed(32'sh0) : $signed(_GEN_4870); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4872 = 6'h3a == _T_3 ? $signed(32'sh0) : $signed(_GEN_4871); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4873 = 6'h3b == _T_3 ? $signed(32'sh0) : $signed(_GEN_4872); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4874 = 6'h3c == _T_3 ? $signed(regsB_3_re) : $signed(_GEN_4873); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4875 = 6'h3d == _T_3 ? $signed(regsB_13_re) : $signed(_GEN_4874); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4876 = 6'h3e == _T_3 ? $signed(regsB_23_re) : $signed(_GEN_4875); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4877 = 6'h3f == _T_3 ? $signed(regsB_33_re) : $signed(_GEN_4876); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4878 = 7'h40 == _GEN_8445 ? $signed(regsB_43_re) : $signed(_GEN_4877); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4879 = 7'h41 == _GEN_8445 ? $signed(regsB_53_re) : $signed(_GEN_4878); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4880 = 7'h42 == _GEN_8445 ? $signed(regsB_63_re) : $signed(_GEN_4879); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4881 = 7'h43 == _GEN_8445 ? $signed(regsB_73_re) : $signed(_GEN_4880); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4882 = 7'h44 == _GEN_8445 ? $signed(regsB_83_re) : $signed(_GEN_4881); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4883 = 7'h45 == _GEN_8445 ? $signed(regsB_93_re) : $signed(_GEN_4882); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4884 = 7'h46 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4883); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4885 = 7'h47 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4884); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4886 = 7'h48 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4885); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4887 = 7'h49 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4886); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4888 = 7'h4a == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4887); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4889 = 7'h4b == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4888); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4890 = 7'h4c == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4889); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4891 = 7'h4d == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4890); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4892 = 7'h4e == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4891); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4893 = 7'h4f == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4892); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4894 = 7'h50 == _GEN_8445 ? $signed(regsB_4_re) : $signed(_GEN_4893); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4895 = 7'h51 == _GEN_8445 ? $signed(regsB_14_re) : $signed(_GEN_4894); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4896 = 7'h52 == _GEN_8445 ? $signed(regsB_24_re) : $signed(_GEN_4895); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4897 = 7'h53 == _GEN_8445 ? $signed(regsB_34_re) : $signed(_GEN_4896); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4898 = 7'h54 == _GEN_8445 ? $signed(regsB_44_re) : $signed(_GEN_4897); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4899 = 7'h55 == _GEN_8445 ? $signed(regsB_54_re) : $signed(_GEN_4898); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4900 = 7'h56 == _GEN_8445 ? $signed(regsB_64_re) : $signed(_GEN_4899); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4901 = 7'h57 == _GEN_8445 ? $signed(regsB_74_re) : $signed(_GEN_4900); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4902 = 7'h58 == _GEN_8445 ? $signed(regsB_84_re) : $signed(_GEN_4901); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4903 = 7'h59 == _GEN_8445 ? $signed(regsB_94_re) : $signed(_GEN_4902); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4904 = 7'h5a == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4903); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4905 = 7'h5b == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4904); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4906 = 7'h5c == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4905); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4907 = 7'h5d == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4906); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4908 = 7'h5e == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4907); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4909 = 7'h5f == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4908); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4910 = 7'h60 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4909); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4911 = 7'h61 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4910); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4912 = 7'h62 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4911); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4913 = 7'h63 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4912); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4914 = 7'h64 == _GEN_8445 ? $signed(regsB_5_re) : $signed(_GEN_4913); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4915 = 7'h65 == _GEN_8445 ? $signed(regsB_15_re) : $signed(_GEN_4914); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4916 = 7'h66 == _GEN_8445 ? $signed(regsB_25_re) : $signed(_GEN_4915); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4917 = 7'h67 == _GEN_8445 ? $signed(regsB_35_re) : $signed(_GEN_4916); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4918 = 7'h68 == _GEN_8445 ? $signed(regsB_45_re) : $signed(_GEN_4917); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4919 = 7'h69 == _GEN_8445 ? $signed(regsB_55_re) : $signed(_GEN_4918); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4920 = 7'h6a == _GEN_8445 ? $signed(regsB_65_re) : $signed(_GEN_4919); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4921 = 7'h6b == _GEN_8445 ? $signed(regsB_75_re) : $signed(_GEN_4920); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4922 = 7'h6c == _GEN_8445 ? $signed(regsB_85_re) : $signed(_GEN_4921); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4923 = 7'h6d == _GEN_8445 ? $signed(regsB_95_re) : $signed(_GEN_4922); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4924 = 7'h6e == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4923); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4925 = 7'h6f == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4924); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4926 = 7'h70 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4925); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4927 = 7'h71 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4926); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4928 = 7'h72 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4927); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4929 = 7'h73 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4928); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4930 = 7'h74 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4929); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4931 = 7'h75 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4930); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4932 = 7'h76 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4931); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4933 = 7'h77 == _GEN_8445 ? $signed(32'sh0) : $signed(_GEN_4932); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4934 = 7'h78 == _GEN_8445 ? $signed(regsB_6_re) : $signed(_GEN_4933); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4935 = 7'h79 == _GEN_8445 ? $signed(regsB_16_re) : $signed(_GEN_4934); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4936 = 7'h7a == _GEN_8445 ? $signed(regsB_26_re) : $signed(_GEN_4935); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4937 = 7'h7b == _GEN_8445 ? $signed(regsB_36_re) : $signed(_GEN_4936); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4938 = 7'h7c == _GEN_8445 ? $signed(regsB_46_re) : $signed(_GEN_4937); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4939 = 7'h7d == _GEN_8445 ? $signed(regsB_56_re) : $signed(_GEN_4938); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4940 = 7'h7e == _GEN_8445 ? $signed(regsB_66_re) : $signed(_GEN_4939); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4941 = 7'h7f == _GEN_8445 ? $signed(regsB_76_re) : $signed(_GEN_4940); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4942 = 8'h80 == _GEN_8509 ? $signed(regsB_86_re) : $signed(_GEN_4941); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4943 = 8'h81 == _GEN_8509 ? $signed(regsB_96_re) : $signed(_GEN_4942); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4944 = 8'h82 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4943); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4945 = 8'h83 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4944); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4946 = 8'h84 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4945); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4947 = 8'h85 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4946); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4948 = 8'h86 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4947); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4949 = 8'h87 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4948); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4950 = 8'h88 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4949); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4951 = 8'h89 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4950); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4952 = 8'h8a == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4951); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4953 = 8'h8b == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4952); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4954 = 8'h8c == _GEN_8509 ? $signed(regsB_7_re) : $signed(_GEN_4953); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4955 = 8'h8d == _GEN_8509 ? $signed(regsB_17_re) : $signed(_GEN_4954); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4956 = 8'h8e == _GEN_8509 ? $signed(regsB_27_re) : $signed(_GEN_4955); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4957 = 8'h8f == _GEN_8509 ? $signed(regsB_37_re) : $signed(_GEN_4956); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4958 = 8'h90 == _GEN_8509 ? $signed(regsB_47_re) : $signed(_GEN_4957); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4959 = 8'h91 == _GEN_8509 ? $signed(regsB_57_re) : $signed(_GEN_4958); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4960 = 8'h92 == _GEN_8509 ? $signed(regsB_67_re) : $signed(_GEN_4959); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4961 = 8'h93 == _GEN_8509 ? $signed(regsB_77_re) : $signed(_GEN_4960); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4962 = 8'h94 == _GEN_8509 ? $signed(regsB_87_re) : $signed(_GEN_4961); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4963 = 8'h95 == _GEN_8509 ? $signed(regsB_97_re) : $signed(_GEN_4962); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4964 = 8'h96 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4963); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4965 = 8'h97 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4964); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4966 = 8'h98 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4965); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4967 = 8'h99 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4966); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4968 = 8'h9a == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4967); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4969 = 8'h9b == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4968); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4970 = 8'h9c == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4969); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4971 = 8'h9d == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4970); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4972 = 8'h9e == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4971); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4973 = 8'h9f == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4972); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4974 = 8'ha0 == _GEN_8509 ? $signed(regsB_8_re) : $signed(_GEN_4973); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4975 = 8'ha1 == _GEN_8509 ? $signed(regsB_18_re) : $signed(_GEN_4974); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4976 = 8'ha2 == _GEN_8509 ? $signed(regsB_28_re) : $signed(_GEN_4975); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4977 = 8'ha3 == _GEN_8509 ? $signed(regsB_38_re) : $signed(_GEN_4976); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4978 = 8'ha4 == _GEN_8509 ? $signed(regsB_48_re) : $signed(_GEN_4977); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4979 = 8'ha5 == _GEN_8509 ? $signed(regsB_58_re) : $signed(_GEN_4978); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4980 = 8'ha6 == _GEN_8509 ? $signed(regsB_68_re) : $signed(_GEN_4979); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4981 = 8'ha7 == _GEN_8509 ? $signed(regsB_78_re) : $signed(_GEN_4980); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4982 = 8'ha8 == _GEN_8509 ? $signed(regsB_88_re) : $signed(_GEN_4981); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4983 = 8'ha9 == _GEN_8509 ? $signed(regsB_98_re) : $signed(_GEN_4982); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4984 = 8'haa == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4983); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4985 = 8'hab == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4984); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4986 = 8'hac == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4985); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4987 = 8'had == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4986); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4988 = 8'hae == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4987); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4989 = 8'haf == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4988); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4990 = 8'hb0 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4989); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4991 = 8'hb1 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4990); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4992 = 8'hb2 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4991); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4993 = 8'hb3 == _GEN_8509 ? $signed(32'sh0) : $signed(_GEN_4992); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4994 = 8'hb4 == _GEN_8509 ? $signed(regsB_9_re) : $signed(_GEN_4993); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4995 = 8'hb5 == _GEN_8509 ? $signed(regsB_19_re) : $signed(_GEN_4994); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4996 = 8'hb6 == _GEN_8509 ? $signed(regsB_29_re) : $signed(_GEN_4995); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4997 = 8'hb7 == _GEN_8509 ? $signed(regsB_39_re) : $signed(_GEN_4996); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4998 = 8'hb8 == _GEN_8509 ? $signed(regsB_49_re) : $signed(_GEN_4997); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_4999 = 8'hb9 == _GEN_8509 ? $signed(regsB_59_re) : $signed(_GEN_4998); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5000 = 8'hba == _GEN_8509 ? $signed(regsB_69_re) : $signed(_GEN_4999); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5001 = 8'hbb == _GEN_8509 ? $signed(regsB_79_re) : $signed(_GEN_5000); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5002 = 8'hbc == _GEN_8509 ? $signed(regsB_89_re) : $signed(_GEN_5001); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5003 = 8'hbd == _GEN_8509 ? $signed(regsB_99_re) : $signed(_GEN_5002); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5005 = 6'h1 == _T_6 ? $signed(regsB_10_im) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5006 = 6'h2 == _T_6 ? $signed(regsB_20_im) : $signed(_GEN_5005); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5007 = 6'h3 == _T_6 ? $signed(regsB_30_im) : $signed(_GEN_5006); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5008 = 6'h4 == _T_6 ? $signed(regsB_40_im) : $signed(_GEN_5007); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5009 = 6'h5 == _T_6 ? $signed(regsB_50_im) : $signed(_GEN_5008); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5010 = 6'h6 == _T_6 ? $signed(regsB_60_im) : $signed(_GEN_5009); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5011 = 6'h7 == _T_6 ? $signed(regsB_70_im) : $signed(_GEN_5010); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5012 = 6'h8 == _T_6 ? $signed(regsB_80_im) : $signed(_GEN_5011); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5013 = 6'h9 == _T_6 ? $signed(regsB_90_im) : $signed(_GEN_5012); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5014 = 6'ha == _T_6 ? $signed(32'sh0) : $signed(_GEN_5013); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5015 = 6'hb == _T_6 ? $signed(32'sh0) : $signed(_GEN_5014); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5016 = 6'hc == _T_6 ? $signed(32'sh0) : $signed(_GEN_5015); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5017 = 6'hd == _T_6 ? $signed(32'sh0) : $signed(_GEN_5016); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5018 = 6'he == _T_6 ? $signed(32'sh0) : $signed(_GEN_5017); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5019 = 6'hf == _T_6 ? $signed(32'sh0) : $signed(_GEN_5018); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5020 = 6'h10 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5019); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5021 = 6'h11 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5020); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5022 = 6'h12 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5021); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5023 = 6'h13 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5022); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5024 = 6'h14 == _T_6 ? $signed(regsB_1_im) : $signed(_GEN_5023); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5025 = 6'h15 == _T_6 ? $signed(regsB_11_im) : $signed(_GEN_5024); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5026 = 6'h16 == _T_6 ? $signed(regsB_21_im) : $signed(_GEN_5025); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5027 = 6'h17 == _T_6 ? $signed(regsB_31_im) : $signed(_GEN_5026); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5028 = 6'h18 == _T_6 ? $signed(regsB_41_im) : $signed(_GEN_5027); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5029 = 6'h19 == _T_6 ? $signed(regsB_51_im) : $signed(_GEN_5028); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5030 = 6'h1a == _T_6 ? $signed(regsB_61_im) : $signed(_GEN_5029); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5031 = 6'h1b == _T_6 ? $signed(regsB_71_im) : $signed(_GEN_5030); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5032 = 6'h1c == _T_6 ? $signed(regsB_81_im) : $signed(_GEN_5031); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5033 = 6'h1d == _T_6 ? $signed(regsB_91_im) : $signed(_GEN_5032); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5034 = 6'h1e == _T_6 ? $signed(32'sh0) : $signed(_GEN_5033); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5035 = 6'h1f == _T_6 ? $signed(32'sh0) : $signed(_GEN_5034); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5036 = 6'h20 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5035); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5037 = 6'h21 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5036); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5038 = 6'h22 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5037); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5039 = 6'h23 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5038); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5040 = 6'h24 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5039); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5041 = 6'h25 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5040); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5042 = 6'h26 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5041); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5043 = 6'h27 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5042); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5044 = 6'h28 == _T_6 ? $signed(regsB_2_im) : $signed(_GEN_5043); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5045 = 6'h29 == _T_6 ? $signed(regsB_12_im) : $signed(_GEN_5044); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5046 = 6'h2a == _T_6 ? $signed(regsB_22_im) : $signed(_GEN_5045); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5047 = 6'h2b == _T_6 ? $signed(regsB_32_im) : $signed(_GEN_5046); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5048 = 6'h2c == _T_6 ? $signed(regsB_42_im) : $signed(_GEN_5047); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5049 = 6'h2d == _T_6 ? $signed(regsB_52_im) : $signed(_GEN_5048); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5050 = 6'h2e == _T_6 ? $signed(regsB_62_im) : $signed(_GEN_5049); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5051 = 6'h2f == _T_6 ? $signed(regsB_72_im) : $signed(_GEN_5050); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5052 = 6'h30 == _T_6 ? $signed(regsB_82_im) : $signed(_GEN_5051); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5053 = 6'h31 == _T_6 ? $signed(regsB_92_im) : $signed(_GEN_5052); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5054 = 6'h32 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5053); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5055 = 6'h33 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5054); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5056 = 6'h34 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5055); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5057 = 6'h35 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5056); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5058 = 6'h36 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5057); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5059 = 6'h37 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5058); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5060 = 6'h38 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5059); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5061 = 6'h39 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5060); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5062 = 6'h3a == _T_6 ? $signed(32'sh0) : $signed(_GEN_5061); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5063 = 6'h3b == _T_6 ? $signed(32'sh0) : $signed(_GEN_5062); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5064 = 6'h3c == _T_6 ? $signed(regsB_3_im) : $signed(_GEN_5063); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5065 = 6'h3d == _T_6 ? $signed(regsB_13_im) : $signed(_GEN_5064); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5066 = 6'h3e == _T_6 ? $signed(regsB_23_im) : $signed(_GEN_5065); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5067 = 6'h3f == _T_6 ? $signed(regsB_33_im) : $signed(_GEN_5066); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5068 = 7'h40 == _GEN_8697 ? $signed(regsB_43_im) : $signed(_GEN_5067); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5069 = 7'h41 == _GEN_8697 ? $signed(regsB_53_im) : $signed(_GEN_5068); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5070 = 7'h42 == _GEN_8697 ? $signed(regsB_63_im) : $signed(_GEN_5069); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5071 = 7'h43 == _GEN_8697 ? $signed(regsB_73_im) : $signed(_GEN_5070); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5072 = 7'h44 == _GEN_8697 ? $signed(regsB_83_im) : $signed(_GEN_5071); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5073 = 7'h45 == _GEN_8697 ? $signed(regsB_93_im) : $signed(_GEN_5072); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5074 = 7'h46 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5073); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5075 = 7'h47 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5074); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5076 = 7'h48 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5075); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5077 = 7'h49 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5076); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5078 = 7'h4a == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5077); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5079 = 7'h4b == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5078); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5080 = 7'h4c == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5079); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5081 = 7'h4d == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5080); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5082 = 7'h4e == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5081); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5083 = 7'h4f == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5082); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5084 = 7'h50 == _GEN_8697 ? $signed(regsB_4_im) : $signed(_GEN_5083); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5085 = 7'h51 == _GEN_8697 ? $signed(regsB_14_im) : $signed(_GEN_5084); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5086 = 7'h52 == _GEN_8697 ? $signed(regsB_24_im) : $signed(_GEN_5085); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5087 = 7'h53 == _GEN_8697 ? $signed(regsB_34_im) : $signed(_GEN_5086); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5088 = 7'h54 == _GEN_8697 ? $signed(regsB_44_im) : $signed(_GEN_5087); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5089 = 7'h55 == _GEN_8697 ? $signed(regsB_54_im) : $signed(_GEN_5088); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5090 = 7'h56 == _GEN_8697 ? $signed(regsB_64_im) : $signed(_GEN_5089); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5091 = 7'h57 == _GEN_8697 ? $signed(regsB_74_im) : $signed(_GEN_5090); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5092 = 7'h58 == _GEN_8697 ? $signed(regsB_84_im) : $signed(_GEN_5091); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5093 = 7'h59 == _GEN_8697 ? $signed(regsB_94_im) : $signed(_GEN_5092); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5094 = 7'h5a == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5093); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5095 = 7'h5b == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5094); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5096 = 7'h5c == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5095); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5097 = 7'h5d == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5096); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5098 = 7'h5e == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5097); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5099 = 7'h5f == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5098); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5100 = 7'h60 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5099); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5101 = 7'h61 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5100); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5102 = 7'h62 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5101); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5103 = 7'h63 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5102); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5104 = 7'h64 == _GEN_8697 ? $signed(regsB_5_im) : $signed(_GEN_5103); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5105 = 7'h65 == _GEN_8697 ? $signed(regsB_15_im) : $signed(_GEN_5104); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5106 = 7'h66 == _GEN_8697 ? $signed(regsB_25_im) : $signed(_GEN_5105); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5107 = 7'h67 == _GEN_8697 ? $signed(regsB_35_im) : $signed(_GEN_5106); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5108 = 7'h68 == _GEN_8697 ? $signed(regsB_45_im) : $signed(_GEN_5107); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5109 = 7'h69 == _GEN_8697 ? $signed(regsB_55_im) : $signed(_GEN_5108); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5110 = 7'h6a == _GEN_8697 ? $signed(regsB_65_im) : $signed(_GEN_5109); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5111 = 7'h6b == _GEN_8697 ? $signed(regsB_75_im) : $signed(_GEN_5110); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5112 = 7'h6c == _GEN_8697 ? $signed(regsB_85_im) : $signed(_GEN_5111); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5113 = 7'h6d == _GEN_8697 ? $signed(regsB_95_im) : $signed(_GEN_5112); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5114 = 7'h6e == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5113); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5115 = 7'h6f == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5114); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5116 = 7'h70 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5115); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5117 = 7'h71 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5116); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5118 = 7'h72 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5117); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5119 = 7'h73 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5118); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5120 = 7'h74 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5119); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5121 = 7'h75 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5120); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5122 = 7'h76 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5121); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5123 = 7'h77 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5122); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5124 = 7'h78 == _GEN_8697 ? $signed(regsB_6_im) : $signed(_GEN_5123); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5125 = 7'h79 == _GEN_8697 ? $signed(regsB_16_im) : $signed(_GEN_5124); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5126 = 7'h7a == _GEN_8697 ? $signed(regsB_26_im) : $signed(_GEN_5125); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5127 = 7'h7b == _GEN_8697 ? $signed(regsB_36_im) : $signed(_GEN_5126); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5128 = 7'h7c == _GEN_8697 ? $signed(regsB_46_im) : $signed(_GEN_5127); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5129 = 7'h7d == _GEN_8697 ? $signed(regsB_56_im) : $signed(_GEN_5128); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5130 = 7'h7e == _GEN_8697 ? $signed(regsB_66_im) : $signed(_GEN_5129); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5131 = 7'h7f == _GEN_8697 ? $signed(regsB_76_im) : $signed(_GEN_5130); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5132 = 8'h80 == _GEN_8761 ? $signed(regsB_86_im) : $signed(_GEN_5131); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5133 = 8'h81 == _GEN_8761 ? $signed(regsB_96_im) : $signed(_GEN_5132); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5134 = 8'h82 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5133); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5135 = 8'h83 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5134); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5136 = 8'h84 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5135); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5137 = 8'h85 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5136); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5138 = 8'h86 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5137); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5139 = 8'h87 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5138); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5140 = 8'h88 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5139); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5141 = 8'h89 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5140); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5142 = 8'h8a == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5141); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5143 = 8'h8b == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5142); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5144 = 8'h8c == _GEN_8761 ? $signed(regsB_7_im) : $signed(_GEN_5143); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5145 = 8'h8d == _GEN_8761 ? $signed(regsB_17_im) : $signed(_GEN_5144); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5146 = 8'h8e == _GEN_8761 ? $signed(regsB_27_im) : $signed(_GEN_5145); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5147 = 8'h8f == _GEN_8761 ? $signed(regsB_37_im) : $signed(_GEN_5146); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5148 = 8'h90 == _GEN_8761 ? $signed(regsB_47_im) : $signed(_GEN_5147); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5149 = 8'h91 == _GEN_8761 ? $signed(regsB_57_im) : $signed(_GEN_5148); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5150 = 8'h92 == _GEN_8761 ? $signed(regsB_67_im) : $signed(_GEN_5149); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5151 = 8'h93 == _GEN_8761 ? $signed(regsB_77_im) : $signed(_GEN_5150); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5152 = 8'h94 == _GEN_8761 ? $signed(regsB_87_im) : $signed(_GEN_5151); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5153 = 8'h95 == _GEN_8761 ? $signed(regsB_97_im) : $signed(_GEN_5152); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5154 = 8'h96 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5153); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5155 = 8'h97 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5154); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5156 = 8'h98 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5155); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5157 = 8'h99 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5156); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5158 = 8'h9a == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5157); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5159 = 8'h9b == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5158); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5160 = 8'h9c == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5159); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5161 = 8'h9d == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5160); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5162 = 8'h9e == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5161); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5163 = 8'h9f == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5162); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5164 = 8'ha0 == _GEN_8761 ? $signed(regsB_8_im) : $signed(_GEN_5163); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5165 = 8'ha1 == _GEN_8761 ? $signed(regsB_18_im) : $signed(_GEN_5164); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5166 = 8'ha2 == _GEN_8761 ? $signed(regsB_28_im) : $signed(_GEN_5165); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5167 = 8'ha3 == _GEN_8761 ? $signed(regsB_38_im) : $signed(_GEN_5166); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5168 = 8'ha4 == _GEN_8761 ? $signed(regsB_48_im) : $signed(_GEN_5167); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5169 = 8'ha5 == _GEN_8761 ? $signed(regsB_58_im) : $signed(_GEN_5168); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5170 = 8'ha6 == _GEN_8761 ? $signed(regsB_68_im) : $signed(_GEN_5169); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5171 = 8'ha7 == _GEN_8761 ? $signed(regsB_78_im) : $signed(_GEN_5170); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5172 = 8'ha8 == _GEN_8761 ? $signed(regsB_88_im) : $signed(_GEN_5171); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5173 = 8'ha9 == _GEN_8761 ? $signed(regsB_98_im) : $signed(_GEN_5172); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5174 = 8'haa == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5173); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5175 = 8'hab == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5174); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5176 = 8'hac == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5175); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5177 = 8'had == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5176); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5178 = 8'hae == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5177); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5179 = 8'haf == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5178); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5180 = 8'hb0 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5179); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5181 = 8'hb1 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5180); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5182 = 8'hb2 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5181); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5183 = 8'hb3 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5182); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5184 = 8'hb4 == _GEN_8761 ? $signed(regsB_9_im) : $signed(_GEN_5183); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5185 = 8'hb5 == _GEN_8761 ? $signed(regsB_19_im) : $signed(_GEN_5184); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5186 = 8'hb6 == _GEN_8761 ? $signed(regsB_29_im) : $signed(_GEN_5185); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5187 = 8'hb7 == _GEN_8761 ? $signed(regsB_39_im) : $signed(_GEN_5186); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5188 = 8'hb8 == _GEN_8761 ? $signed(regsB_49_im) : $signed(_GEN_5187); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5189 = 8'hb9 == _GEN_8761 ? $signed(regsB_59_im) : $signed(_GEN_5188); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5190 = 8'hba == _GEN_8761 ? $signed(regsB_69_im) : $signed(_GEN_5189); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5191 = 8'hbb == _GEN_8761 ? $signed(regsB_79_im) : $signed(_GEN_5190); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5192 = 8'hbc == _GEN_8761 ? $signed(regsB_89_im) : $signed(_GEN_5191); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5193 = 8'hbd == _GEN_8761 ? $signed(regsB_99_im) : $signed(_GEN_5192); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5195 = 6'h1 == _T_6 ? $signed(regsB_10_re) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5196 = 6'h2 == _T_6 ? $signed(regsB_20_re) : $signed(_GEN_5195); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5197 = 6'h3 == _T_6 ? $signed(regsB_30_re) : $signed(_GEN_5196); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5198 = 6'h4 == _T_6 ? $signed(regsB_40_re) : $signed(_GEN_5197); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5199 = 6'h5 == _T_6 ? $signed(regsB_50_re) : $signed(_GEN_5198); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5200 = 6'h6 == _T_6 ? $signed(regsB_60_re) : $signed(_GEN_5199); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5201 = 6'h7 == _T_6 ? $signed(regsB_70_re) : $signed(_GEN_5200); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5202 = 6'h8 == _T_6 ? $signed(regsB_80_re) : $signed(_GEN_5201); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5203 = 6'h9 == _T_6 ? $signed(regsB_90_re) : $signed(_GEN_5202); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5204 = 6'ha == _T_6 ? $signed(32'sh0) : $signed(_GEN_5203); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5205 = 6'hb == _T_6 ? $signed(32'sh0) : $signed(_GEN_5204); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5206 = 6'hc == _T_6 ? $signed(32'sh0) : $signed(_GEN_5205); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5207 = 6'hd == _T_6 ? $signed(32'sh0) : $signed(_GEN_5206); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5208 = 6'he == _T_6 ? $signed(32'sh0) : $signed(_GEN_5207); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5209 = 6'hf == _T_6 ? $signed(32'sh0) : $signed(_GEN_5208); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5210 = 6'h10 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5209); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5211 = 6'h11 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5210); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5212 = 6'h12 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5211); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5213 = 6'h13 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5212); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5214 = 6'h14 == _T_6 ? $signed(regsB_1_re) : $signed(_GEN_5213); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5215 = 6'h15 == _T_6 ? $signed(regsB_11_re) : $signed(_GEN_5214); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5216 = 6'h16 == _T_6 ? $signed(regsB_21_re) : $signed(_GEN_5215); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5217 = 6'h17 == _T_6 ? $signed(regsB_31_re) : $signed(_GEN_5216); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5218 = 6'h18 == _T_6 ? $signed(regsB_41_re) : $signed(_GEN_5217); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5219 = 6'h19 == _T_6 ? $signed(regsB_51_re) : $signed(_GEN_5218); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5220 = 6'h1a == _T_6 ? $signed(regsB_61_re) : $signed(_GEN_5219); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5221 = 6'h1b == _T_6 ? $signed(regsB_71_re) : $signed(_GEN_5220); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5222 = 6'h1c == _T_6 ? $signed(regsB_81_re) : $signed(_GEN_5221); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5223 = 6'h1d == _T_6 ? $signed(regsB_91_re) : $signed(_GEN_5222); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5224 = 6'h1e == _T_6 ? $signed(32'sh0) : $signed(_GEN_5223); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5225 = 6'h1f == _T_6 ? $signed(32'sh0) : $signed(_GEN_5224); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5226 = 6'h20 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5225); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5227 = 6'h21 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5226); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5228 = 6'h22 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5227); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5229 = 6'h23 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5228); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5230 = 6'h24 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5229); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5231 = 6'h25 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5230); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5232 = 6'h26 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5231); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5233 = 6'h27 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5232); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5234 = 6'h28 == _T_6 ? $signed(regsB_2_re) : $signed(_GEN_5233); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5235 = 6'h29 == _T_6 ? $signed(regsB_12_re) : $signed(_GEN_5234); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5236 = 6'h2a == _T_6 ? $signed(regsB_22_re) : $signed(_GEN_5235); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5237 = 6'h2b == _T_6 ? $signed(regsB_32_re) : $signed(_GEN_5236); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5238 = 6'h2c == _T_6 ? $signed(regsB_42_re) : $signed(_GEN_5237); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5239 = 6'h2d == _T_6 ? $signed(regsB_52_re) : $signed(_GEN_5238); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5240 = 6'h2e == _T_6 ? $signed(regsB_62_re) : $signed(_GEN_5239); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5241 = 6'h2f == _T_6 ? $signed(regsB_72_re) : $signed(_GEN_5240); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5242 = 6'h30 == _T_6 ? $signed(regsB_82_re) : $signed(_GEN_5241); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5243 = 6'h31 == _T_6 ? $signed(regsB_92_re) : $signed(_GEN_5242); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5244 = 6'h32 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5243); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5245 = 6'h33 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5244); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5246 = 6'h34 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5245); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5247 = 6'h35 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5246); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5248 = 6'h36 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5247); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5249 = 6'h37 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5248); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5250 = 6'h38 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5249); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5251 = 6'h39 == _T_6 ? $signed(32'sh0) : $signed(_GEN_5250); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5252 = 6'h3a == _T_6 ? $signed(32'sh0) : $signed(_GEN_5251); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5253 = 6'h3b == _T_6 ? $signed(32'sh0) : $signed(_GEN_5252); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5254 = 6'h3c == _T_6 ? $signed(regsB_3_re) : $signed(_GEN_5253); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5255 = 6'h3d == _T_6 ? $signed(regsB_13_re) : $signed(_GEN_5254); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5256 = 6'h3e == _T_6 ? $signed(regsB_23_re) : $signed(_GEN_5255); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5257 = 6'h3f == _T_6 ? $signed(regsB_33_re) : $signed(_GEN_5256); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5258 = 7'h40 == _GEN_8697 ? $signed(regsB_43_re) : $signed(_GEN_5257); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5259 = 7'h41 == _GEN_8697 ? $signed(regsB_53_re) : $signed(_GEN_5258); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5260 = 7'h42 == _GEN_8697 ? $signed(regsB_63_re) : $signed(_GEN_5259); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5261 = 7'h43 == _GEN_8697 ? $signed(regsB_73_re) : $signed(_GEN_5260); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5262 = 7'h44 == _GEN_8697 ? $signed(regsB_83_re) : $signed(_GEN_5261); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5263 = 7'h45 == _GEN_8697 ? $signed(regsB_93_re) : $signed(_GEN_5262); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5264 = 7'h46 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5263); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5265 = 7'h47 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5264); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5266 = 7'h48 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5265); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5267 = 7'h49 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5266); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5268 = 7'h4a == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5267); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5269 = 7'h4b == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5268); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5270 = 7'h4c == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5269); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5271 = 7'h4d == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5270); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5272 = 7'h4e == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5271); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5273 = 7'h4f == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5272); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5274 = 7'h50 == _GEN_8697 ? $signed(regsB_4_re) : $signed(_GEN_5273); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5275 = 7'h51 == _GEN_8697 ? $signed(regsB_14_re) : $signed(_GEN_5274); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5276 = 7'h52 == _GEN_8697 ? $signed(regsB_24_re) : $signed(_GEN_5275); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5277 = 7'h53 == _GEN_8697 ? $signed(regsB_34_re) : $signed(_GEN_5276); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5278 = 7'h54 == _GEN_8697 ? $signed(regsB_44_re) : $signed(_GEN_5277); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5279 = 7'h55 == _GEN_8697 ? $signed(regsB_54_re) : $signed(_GEN_5278); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5280 = 7'h56 == _GEN_8697 ? $signed(regsB_64_re) : $signed(_GEN_5279); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5281 = 7'h57 == _GEN_8697 ? $signed(regsB_74_re) : $signed(_GEN_5280); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5282 = 7'h58 == _GEN_8697 ? $signed(regsB_84_re) : $signed(_GEN_5281); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5283 = 7'h59 == _GEN_8697 ? $signed(regsB_94_re) : $signed(_GEN_5282); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5284 = 7'h5a == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5283); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5285 = 7'h5b == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5284); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5286 = 7'h5c == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5285); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5287 = 7'h5d == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5286); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5288 = 7'h5e == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5287); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5289 = 7'h5f == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5288); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5290 = 7'h60 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5289); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5291 = 7'h61 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5290); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5292 = 7'h62 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5291); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5293 = 7'h63 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5292); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5294 = 7'h64 == _GEN_8697 ? $signed(regsB_5_re) : $signed(_GEN_5293); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5295 = 7'h65 == _GEN_8697 ? $signed(regsB_15_re) : $signed(_GEN_5294); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5296 = 7'h66 == _GEN_8697 ? $signed(regsB_25_re) : $signed(_GEN_5295); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5297 = 7'h67 == _GEN_8697 ? $signed(regsB_35_re) : $signed(_GEN_5296); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5298 = 7'h68 == _GEN_8697 ? $signed(regsB_45_re) : $signed(_GEN_5297); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5299 = 7'h69 == _GEN_8697 ? $signed(regsB_55_re) : $signed(_GEN_5298); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5300 = 7'h6a == _GEN_8697 ? $signed(regsB_65_re) : $signed(_GEN_5299); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5301 = 7'h6b == _GEN_8697 ? $signed(regsB_75_re) : $signed(_GEN_5300); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5302 = 7'h6c == _GEN_8697 ? $signed(regsB_85_re) : $signed(_GEN_5301); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5303 = 7'h6d == _GEN_8697 ? $signed(regsB_95_re) : $signed(_GEN_5302); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5304 = 7'h6e == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5303); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5305 = 7'h6f == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5304); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5306 = 7'h70 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5305); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5307 = 7'h71 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5306); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5308 = 7'h72 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5307); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5309 = 7'h73 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5308); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5310 = 7'h74 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5309); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5311 = 7'h75 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5310); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5312 = 7'h76 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5311); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5313 = 7'h77 == _GEN_8697 ? $signed(32'sh0) : $signed(_GEN_5312); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5314 = 7'h78 == _GEN_8697 ? $signed(regsB_6_re) : $signed(_GEN_5313); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5315 = 7'h79 == _GEN_8697 ? $signed(regsB_16_re) : $signed(_GEN_5314); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5316 = 7'h7a == _GEN_8697 ? $signed(regsB_26_re) : $signed(_GEN_5315); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5317 = 7'h7b == _GEN_8697 ? $signed(regsB_36_re) : $signed(_GEN_5316); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5318 = 7'h7c == _GEN_8697 ? $signed(regsB_46_re) : $signed(_GEN_5317); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5319 = 7'h7d == _GEN_8697 ? $signed(regsB_56_re) : $signed(_GEN_5318); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5320 = 7'h7e == _GEN_8697 ? $signed(regsB_66_re) : $signed(_GEN_5319); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5321 = 7'h7f == _GEN_8697 ? $signed(regsB_76_re) : $signed(_GEN_5320); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5322 = 8'h80 == _GEN_8761 ? $signed(regsB_86_re) : $signed(_GEN_5321); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5323 = 8'h81 == _GEN_8761 ? $signed(regsB_96_re) : $signed(_GEN_5322); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5324 = 8'h82 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5323); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5325 = 8'h83 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5324); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5326 = 8'h84 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5325); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5327 = 8'h85 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5326); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5328 = 8'h86 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5327); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5329 = 8'h87 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5328); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5330 = 8'h88 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5329); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5331 = 8'h89 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5330); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5332 = 8'h8a == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5331); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5333 = 8'h8b == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5332); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5334 = 8'h8c == _GEN_8761 ? $signed(regsB_7_re) : $signed(_GEN_5333); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5335 = 8'h8d == _GEN_8761 ? $signed(regsB_17_re) : $signed(_GEN_5334); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5336 = 8'h8e == _GEN_8761 ? $signed(regsB_27_re) : $signed(_GEN_5335); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5337 = 8'h8f == _GEN_8761 ? $signed(regsB_37_re) : $signed(_GEN_5336); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5338 = 8'h90 == _GEN_8761 ? $signed(regsB_47_re) : $signed(_GEN_5337); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5339 = 8'h91 == _GEN_8761 ? $signed(regsB_57_re) : $signed(_GEN_5338); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5340 = 8'h92 == _GEN_8761 ? $signed(regsB_67_re) : $signed(_GEN_5339); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5341 = 8'h93 == _GEN_8761 ? $signed(regsB_77_re) : $signed(_GEN_5340); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5342 = 8'h94 == _GEN_8761 ? $signed(regsB_87_re) : $signed(_GEN_5341); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5343 = 8'h95 == _GEN_8761 ? $signed(regsB_97_re) : $signed(_GEN_5342); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5344 = 8'h96 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5343); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5345 = 8'h97 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5344); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5346 = 8'h98 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5345); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5347 = 8'h99 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5346); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5348 = 8'h9a == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5347); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5349 = 8'h9b == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5348); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5350 = 8'h9c == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5349); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5351 = 8'h9d == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5350); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5352 = 8'h9e == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5351); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5353 = 8'h9f == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5352); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5354 = 8'ha0 == _GEN_8761 ? $signed(regsB_8_re) : $signed(_GEN_5353); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5355 = 8'ha1 == _GEN_8761 ? $signed(regsB_18_re) : $signed(_GEN_5354); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5356 = 8'ha2 == _GEN_8761 ? $signed(regsB_28_re) : $signed(_GEN_5355); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5357 = 8'ha3 == _GEN_8761 ? $signed(regsB_38_re) : $signed(_GEN_5356); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5358 = 8'ha4 == _GEN_8761 ? $signed(regsB_48_re) : $signed(_GEN_5357); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5359 = 8'ha5 == _GEN_8761 ? $signed(regsB_58_re) : $signed(_GEN_5358); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5360 = 8'ha6 == _GEN_8761 ? $signed(regsB_68_re) : $signed(_GEN_5359); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5361 = 8'ha7 == _GEN_8761 ? $signed(regsB_78_re) : $signed(_GEN_5360); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5362 = 8'ha8 == _GEN_8761 ? $signed(regsB_88_re) : $signed(_GEN_5361); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5363 = 8'ha9 == _GEN_8761 ? $signed(regsB_98_re) : $signed(_GEN_5362); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5364 = 8'haa == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5363); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5365 = 8'hab == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5364); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5366 = 8'hac == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5365); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5367 = 8'had == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5366); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5368 = 8'hae == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5367); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5369 = 8'haf == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5368); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5370 = 8'hb0 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5369); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5371 = 8'hb1 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5370); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5372 = 8'hb2 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5371); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5373 = 8'hb3 == _GEN_8761 ? $signed(32'sh0) : $signed(_GEN_5372); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5374 = 8'hb4 == _GEN_8761 ? $signed(regsB_9_re) : $signed(_GEN_5373); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5375 = 8'hb5 == _GEN_8761 ? $signed(regsB_19_re) : $signed(_GEN_5374); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5376 = 8'hb6 == _GEN_8761 ? $signed(regsB_29_re) : $signed(_GEN_5375); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5377 = 8'hb7 == _GEN_8761 ? $signed(regsB_39_re) : $signed(_GEN_5376); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5378 = 8'hb8 == _GEN_8761 ? $signed(regsB_49_re) : $signed(_GEN_5377); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5379 = 8'hb9 == _GEN_8761 ? $signed(regsB_59_re) : $signed(_GEN_5378); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5380 = 8'hba == _GEN_8761 ? $signed(regsB_69_re) : $signed(_GEN_5379); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5381 = 8'hbb == _GEN_8761 ? $signed(regsB_79_re) : $signed(_GEN_5380); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5382 = 8'hbc == _GEN_8761 ? $signed(regsB_89_re) : $signed(_GEN_5381); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5383 = 8'hbd == _GEN_8761 ? $signed(regsB_99_re) : $signed(_GEN_5382); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5385 = 7'h1 == _T_9 ? $signed(regsB_10_im) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5386 = 7'h2 == _T_9 ? $signed(regsB_20_im) : $signed(_GEN_5385); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5387 = 7'h3 == _T_9 ? $signed(regsB_30_im) : $signed(_GEN_5386); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5388 = 7'h4 == _T_9 ? $signed(regsB_40_im) : $signed(_GEN_5387); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5389 = 7'h5 == _T_9 ? $signed(regsB_50_im) : $signed(_GEN_5388); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5390 = 7'h6 == _T_9 ? $signed(regsB_60_im) : $signed(_GEN_5389); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5391 = 7'h7 == _T_9 ? $signed(regsB_70_im) : $signed(_GEN_5390); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5392 = 7'h8 == _T_9 ? $signed(regsB_80_im) : $signed(_GEN_5391); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5393 = 7'h9 == _T_9 ? $signed(regsB_90_im) : $signed(_GEN_5392); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5394 = 7'ha == _T_9 ? $signed(32'sh0) : $signed(_GEN_5393); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5395 = 7'hb == _T_9 ? $signed(32'sh0) : $signed(_GEN_5394); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5396 = 7'hc == _T_9 ? $signed(32'sh0) : $signed(_GEN_5395); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5397 = 7'hd == _T_9 ? $signed(32'sh0) : $signed(_GEN_5396); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5398 = 7'he == _T_9 ? $signed(32'sh0) : $signed(_GEN_5397); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5399 = 7'hf == _T_9 ? $signed(32'sh0) : $signed(_GEN_5398); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5400 = 7'h10 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5399); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5401 = 7'h11 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5400); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5402 = 7'h12 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5401); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5403 = 7'h13 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5402); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5404 = 7'h14 == _T_9 ? $signed(regsB_1_im) : $signed(_GEN_5403); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5405 = 7'h15 == _T_9 ? $signed(regsB_11_im) : $signed(_GEN_5404); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5406 = 7'h16 == _T_9 ? $signed(regsB_21_im) : $signed(_GEN_5405); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5407 = 7'h17 == _T_9 ? $signed(regsB_31_im) : $signed(_GEN_5406); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5408 = 7'h18 == _T_9 ? $signed(regsB_41_im) : $signed(_GEN_5407); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5409 = 7'h19 == _T_9 ? $signed(regsB_51_im) : $signed(_GEN_5408); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5410 = 7'h1a == _T_9 ? $signed(regsB_61_im) : $signed(_GEN_5409); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5411 = 7'h1b == _T_9 ? $signed(regsB_71_im) : $signed(_GEN_5410); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5412 = 7'h1c == _T_9 ? $signed(regsB_81_im) : $signed(_GEN_5411); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5413 = 7'h1d == _T_9 ? $signed(regsB_91_im) : $signed(_GEN_5412); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5414 = 7'h1e == _T_9 ? $signed(32'sh0) : $signed(_GEN_5413); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5415 = 7'h1f == _T_9 ? $signed(32'sh0) : $signed(_GEN_5414); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5416 = 7'h20 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5415); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5417 = 7'h21 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5416); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5418 = 7'h22 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5417); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5419 = 7'h23 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5418); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5420 = 7'h24 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5419); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5421 = 7'h25 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5420); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5422 = 7'h26 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5421); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5423 = 7'h27 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5422); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5424 = 7'h28 == _T_9 ? $signed(regsB_2_im) : $signed(_GEN_5423); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5425 = 7'h29 == _T_9 ? $signed(regsB_12_im) : $signed(_GEN_5424); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5426 = 7'h2a == _T_9 ? $signed(regsB_22_im) : $signed(_GEN_5425); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5427 = 7'h2b == _T_9 ? $signed(regsB_32_im) : $signed(_GEN_5426); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5428 = 7'h2c == _T_9 ? $signed(regsB_42_im) : $signed(_GEN_5427); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5429 = 7'h2d == _T_9 ? $signed(regsB_52_im) : $signed(_GEN_5428); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5430 = 7'h2e == _T_9 ? $signed(regsB_62_im) : $signed(_GEN_5429); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5431 = 7'h2f == _T_9 ? $signed(regsB_72_im) : $signed(_GEN_5430); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5432 = 7'h30 == _T_9 ? $signed(regsB_82_im) : $signed(_GEN_5431); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5433 = 7'h31 == _T_9 ? $signed(regsB_92_im) : $signed(_GEN_5432); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5434 = 7'h32 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5433); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5435 = 7'h33 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5434); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5436 = 7'h34 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5435); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5437 = 7'h35 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5436); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5438 = 7'h36 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5437); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5439 = 7'h37 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5438); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5440 = 7'h38 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5439); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5441 = 7'h39 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5440); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5442 = 7'h3a == _T_9 ? $signed(32'sh0) : $signed(_GEN_5441); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5443 = 7'h3b == _T_9 ? $signed(32'sh0) : $signed(_GEN_5442); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5444 = 7'h3c == _T_9 ? $signed(regsB_3_im) : $signed(_GEN_5443); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5445 = 7'h3d == _T_9 ? $signed(regsB_13_im) : $signed(_GEN_5444); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5446 = 7'h3e == _T_9 ? $signed(regsB_23_im) : $signed(_GEN_5445); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5447 = 7'h3f == _T_9 ? $signed(regsB_33_im) : $signed(_GEN_5446); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5448 = 7'h40 == _T_9 ? $signed(regsB_43_im) : $signed(_GEN_5447); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5449 = 7'h41 == _T_9 ? $signed(regsB_53_im) : $signed(_GEN_5448); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5450 = 7'h42 == _T_9 ? $signed(regsB_63_im) : $signed(_GEN_5449); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5451 = 7'h43 == _T_9 ? $signed(regsB_73_im) : $signed(_GEN_5450); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5452 = 7'h44 == _T_9 ? $signed(regsB_83_im) : $signed(_GEN_5451); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5453 = 7'h45 == _T_9 ? $signed(regsB_93_im) : $signed(_GEN_5452); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5454 = 7'h46 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5453); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5455 = 7'h47 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5454); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5456 = 7'h48 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5455); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5457 = 7'h49 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5456); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5458 = 7'h4a == _T_9 ? $signed(32'sh0) : $signed(_GEN_5457); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5459 = 7'h4b == _T_9 ? $signed(32'sh0) : $signed(_GEN_5458); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5460 = 7'h4c == _T_9 ? $signed(32'sh0) : $signed(_GEN_5459); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5461 = 7'h4d == _T_9 ? $signed(32'sh0) : $signed(_GEN_5460); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5462 = 7'h4e == _T_9 ? $signed(32'sh0) : $signed(_GEN_5461); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5463 = 7'h4f == _T_9 ? $signed(32'sh0) : $signed(_GEN_5462); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5464 = 7'h50 == _T_9 ? $signed(regsB_4_im) : $signed(_GEN_5463); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5465 = 7'h51 == _T_9 ? $signed(regsB_14_im) : $signed(_GEN_5464); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5466 = 7'h52 == _T_9 ? $signed(regsB_24_im) : $signed(_GEN_5465); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5467 = 7'h53 == _T_9 ? $signed(regsB_34_im) : $signed(_GEN_5466); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5468 = 7'h54 == _T_9 ? $signed(regsB_44_im) : $signed(_GEN_5467); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5469 = 7'h55 == _T_9 ? $signed(regsB_54_im) : $signed(_GEN_5468); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5470 = 7'h56 == _T_9 ? $signed(regsB_64_im) : $signed(_GEN_5469); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5471 = 7'h57 == _T_9 ? $signed(regsB_74_im) : $signed(_GEN_5470); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5472 = 7'h58 == _T_9 ? $signed(regsB_84_im) : $signed(_GEN_5471); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5473 = 7'h59 == _T_9 ? $signed(regsB_94_im) : $signed(_GEN_5472); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5474 = 7'h5a == _T_9 ? $signed(32'sh0) : $signed(_GEN_5473); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5475 = 7'h5b == _T_9 ? $signed(32'sh0) : $signed(_GEN_5474); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5476 = 7'h5c == _T_9 ? $signed(32'sh0) : $signed(_GEN_5475); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5477 = 7'h5d == _T_9 ? $signed(32'sh0) : $signed(_GEN_5476); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5478 = 7'h5e == _T_9 ? $signed(32'sh0) : $signed(_GEN_5477); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5479 = 7'h5f == _T_9 ? $signed(32'sh0) : $signed(_GEN_5478); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5480 = 7'h60 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5479); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5481 = 7'h61 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5480); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5482 = 7'h62 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5481); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5483 = 7'h63 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5482); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5484 = 7'h64 == _T_9 ? $signed(regsB_5_im) : $signed(_GEN_5483); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5485 = 7'h65 == _T_9 ? $signed(regsB_15_im) : $signed(_GEN_5484); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5486 = 7'h66 == _T_9 ? $signed(regsB_25_im) : $signed(_GEN_5485); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5487 = 7'h67 == _T_9 ? $signed(regsB_35_im) : $signed(_GEN_5486); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5488 = 7'h68 == _T_9 ? $signed(regsB_45_im) : $signed(_GEN_5487); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5489 = 7'h69 == _T_9 ? $signed(regsB_55_im) : $signed(_GEN_5488); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5490 = 7'h6a == _T_9 ? $signed(regsB_65_im) : $signed(_GEN_5489); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5491 = 7'h6b == _T_9 ? $signed(regsB_75_im) : $signed(_GEN_5490); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5492 = 7'h6c == _T_9 ? $signed(regsB_85_im) : $signed(_GEN_5491); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5493 = 7'h6d == _T_9 ? $signed(regsB_95_im) : $signed(_GEN_5492); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5494 = 7'h6e == _T_9 ? $signed(32'sh0) : $signed(_GEN_5493); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5495 = 7'h6f == _T_9 ? $signed(32'sh0) : $signed(_GEN_5494); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5496 = 7'h70 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5495); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5497 = 7'h71 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5496); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5498 = 7'h72 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5497); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5499 = 7'h73 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5498); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5500 = 7'h74 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5499); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5501 = 7'h75 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5500); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5502 = 7'h76 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5501); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5503 = 7'h77 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5502); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5504 = 7'h78 == _T_9 ? $signed(regsB_6_im) : $signed(_GEN_5503); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5505 = 7'h79 == _T_9 ? $signed(regsB_16_im) : $signed(_GEN_5504); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5506 = 7'h7a == _T_9 ? $signed(regsB_26_im) : $signed(_GEN_5505); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5507 = 7'h7b == _T_9 ? $signed(regsB_36_im) : $signed(_GEN_5506); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5508 = 7'h7c == _T_9 ? $signed(regsB_46_im) : $signed(_GEN_5507); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5509 = 7'h7d == _T_9 ? $signed(regsB_56_im) : $signed(_GEN_5508); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5510 = 7'h7e == _T_9 ? $signed(regsB_66_im) : $signed(_GEN_5509); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5511 = 7'h7f == _T_9 ? $signed(regsB_76_im) : $signed(_GEN_5510); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5512 = 8'h80 == _GEN_8950 ? $signed(regsB_86_im) : $signed(_GEN_5511); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5513 = 8'h81 == _GEN_8950 ? $signed(regsB_96_im) : $signed(_GEN_5512); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5514 = 8'h82 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5513); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5515 = 8'h83 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5514); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5516 = 8'h84 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5515); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5517 = 8'h85 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5516); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5518 = 8'h86 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5517); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5519 = 8'h87 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5518); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5520 = 8'h88 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5519); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5521 = 8'h89 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5520); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5522 = 8'h8a == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5521); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5523 = 8'h8b == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5522); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5524 = 8'h8c == _GEN_8950 ? $signed(regsB_7_im) : $signed(_GEN_5523); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5525 = 8'h8d == _GEN_8950 ? $signed(regsB_17_im) : $signed(_GEN_5524); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5526 = 8'h8e == _GEN_8950 ? $signed(regsB_27_im) : $signed(_GEN_5525); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5527 = 8'h8f == _GEN_8950 ? $signed(regsB_37_im) : $signed(_GEN_5526); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5528 = 8'h90 == _GEN_8950 ? $signed(regsB_47_im) : $signed(_GEN_5527); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5529 = 8'h91 == _GEN_8950 ? $signed(regsB_57_im) : $signed(_GEN_5528); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5530 = 8'h92 == _GEN_8950 ? $signed(regsB_67_im) : $signed(_GEN_5529); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5531 = 8'h93 == _GEN_8950 ? $signed(regsB_77_im) : $signed(_GEN_5530); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5532 = 8'h94 == _GEN_8950 ? $signed(regsB_87_im) : $signed(_GEN_5531); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5533 = 8'h95 == _GEN_8950 ? $signed(regsB_97_im) : $signed(_GEN_5532); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5534 = 8'h96 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5533); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5535 = 8'h97 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5534); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5536 = 8'h98 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5535); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5537 = 8'h99 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5536); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5538 = 8'h9a == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5537); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5539 = 8'h9b == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5538); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5540 = 8'h9c == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5539); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5541 = 8'h9d == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5540); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5542 = 8'h9e == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5541); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5543 = 8'h9f == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5542); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5544 = 8'ha0 == _GEN_8950 ? $signed(regsB_8_im) : $signed(_GEN_5543); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5545 = 8'ha1 == _GEN_8950 ? $signed(regsB_18_im) : $signed(_GEN_5544); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5546 = 8'ha2 == _GEN_8950 ? $signed(regsB_28_im) : $signed(_GEN_5545); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5547 = 8'ha3 == _GEN_8950 ? $signed(regsB_38_im) : $signed(_GEN_5546); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5548 = 8'ha4 == _GEN_8950 ? $signed(regsB_48_im) : $signed(_GEN_5547); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5549 = 8'ha5 == _GEN_8950 ? $signed(regsB_58_im) : $signed(_GEN_5548); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5550 = 8'ha6 == _GEN_8950 ? $signed(regsB_68_im) : $signed(_GEN_5549); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5551 = 8'ha7 == _GEN_8950 ? $signed(regsB_78_im) : $signed(_GEN_5550); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5552 = 8'ha8 == _GEN_8950 ? $signed(regsB_88_im) : $signed(_GEN_5551); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5553 = 8'ha9 == _GEN_8950 ? $signed(regsB_98_im) : $signed(_GEN_5552); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5554 = 8'haa == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5553); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5555 = 8'hab == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5554); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5556 = 8'hac == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5555); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5557 = 8'had == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5556); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5558 = 8'hae == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5557); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5559 = 8'haf == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5558); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5560 = 8'hb0 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5559); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5561 = 8'hb1 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5560); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5562 = 8'hb2 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5561); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5563 = 8'hb3 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5562); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5564 = 8'hb4 == _GEN_8950 ? $signed(regsB_9_im) : $signed(_GEN_5563); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5565 = 8'hb5 == _GEN_8950 ? $signed(regsB_19_im) : $signed(_GEN_5564); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5566 = 8'hb6 == _GEN_8950 ? $signed(regsB_29_im) : $signed(_GEN_5565); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5567 = 8'hb7 == _GEN_8950 ? $signed(regsB_39_im) : $signed(_GEN_5566); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5568 = 8'hb8 == _GEN_8950 ? $signed(regsB_49_im) : $signed(_GEN_5567); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5569 = 8'hb9 == _GEN_8950 ? $signed(regsB_59_im) : $signed(_GEN_5568); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5570 = 8'hba == _GEN_8950 ? $signed(regsB_69_im) : $signed(_GEN_5569); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5571 = 8'hbb == _GEN_8950 ? $signed(regsB_79_im) : $signed(_GEN_5570); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5572 = 8'hbc == _GEN_8950 ? $signed(regsB_89_im) : $signed(_GEN_5571); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5573 = 8'hbd == _GEN_8950 ? $signed(regsB_99_im) : $signed(_GEN_5572); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5575 = 7'h1 == _T_9 ? $signed(regsB_10_re) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5576 = 7'h2 == _T_9 ? $signed(regsB_20_re) : $signed(_GEN_5575); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5577 = 7'h3 == _T_9 ? $signed(regsB_30_re) : $signed(_GEN_5576); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5578 = 7'h4 == _T_9 ? $signed(regsB_40_re) : $signed(_GEN_5577); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5579 = 7'h5 == _T_9 ? $signed(regsB_50_re) : $signed(_GEN_5578); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5580 = 7'h6 == _T_9 ? $signed(regsB_60_re) : $signed(_GEN_5579); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5581 = 7'h7 == _T_9 ? $signed(regsB_70_re) : $signed(_GEN_5580); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5582 = 7'h8 == _T_9 ? $signed(regsB_80_re) : $signed(_GEN_5581); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5583 = 7'h9 == _T_9 ? $signed(regsB_90_re) : $signed(_GEN_5582); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5584 = 7'ha == _T_9 ? $signed(32'sh0) : $signed(_GEN_5583); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5585 = 7'hb == _T_9 ? $signed(32'sh0) : $signed(_GEN_5584); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5586 = 7'hc == _T_9 ? $signed(32'sh0) : $signed(_GEN_5585); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5587 = 7'hd == _T_9 ? $signed(32'sh0) : $signed(_GEN_5586); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5588 = 7'he == _T_9 ? $signed(32'sh0) : $signed(_GEN_5587); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5589 = 7'hf == _T_9 ? $signed(32'sh0) : $signed(_GEN_5588); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5590 = 7'h10 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5589); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5591 = 7'h11 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5590); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5592 = 7'h12 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5591); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5593 = 7'h13 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5592); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5594 = 7'h14 == _T_9 ? $signed(regsB_1_re) : $signed(_GEN_5593); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5595 = 7'h15 == _T_9 ? $signed(regsB_11_re) : $signed(_GEN_5594); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5596 = 7'h16 == _T_9 ? $signed(regsB_21_re) : $signed(_GEN_5595); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5597 = 7'h17 == _T_9 ? $signed(regsB_31_re) : $signed(_GEN_5596); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5598 = 7'h18 == _T_9 ? $signed(regsB_41_re) : $signed(_GEN_5597); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5599 = 7'h19 == _T_9 ? $signed(regsB_51_re) : $signed(_GEN_5598); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5600 = 7'h1a == _T_9 ? $signed(regsB_61_re) : $signed(_GEN_5599); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5601 = 7'h1b == _T_9 ? $signed(regsB_71_re) : $signed(_GEN_5600); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5602 = 7'h1c == _T_9 ? $signed(regsB_81_re) : $signed(_GEN_5601); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5603 = 7'h1d == _T_9 ? $signed(regsB_91_re) : $signed(_GEN_5602); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5604 = 7'h1e == _T_9 ? $signed(32'sh0) : $signed(_GEN_5603); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5605 = 7'h1f == _T_9 ? $signed(32'sh0) : $signed(_GEN_5604); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5606 = 7'h20 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5605); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5607 = 7'h21 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5606); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5608 = 7'h22 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5607); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5609 = 7'h23 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5608); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5610 = 7'h24 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5609); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5611 = 7'h25 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5610); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5612 = 7'h26 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5611); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5613 = 7'h27 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5612); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5614 = 7'h28 == _T_9 ? $signed(regsB_2_re) : $signed(_GEN_5613); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5615 = 7'h29 == _T_9 ? $signed(regsB_12_re) : $signed(_GEN_5614); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5616 = 7'h2a == _T_9 ? $signed(regsB_22_re) : $signed(_GEN_5615); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5617 = 7'h2b == _T_9 ? $signed(regsB_32_re) : $signed(_GEN_5616); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5618 = 7'h2c == _T_9 ? $signed(regsB_42_re) : $signed(_GEN_5617); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5619 = 7'h2d == _T_9 ? $signed(regsB_52_re) : $signed(_GEN_5618); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5620 = 7'h2e == _T_9 ? $signed(regsB_62_re) : $signed(_GEN_5619); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5621 = 7'h2f == _T_9 ? $signed(regsB_72_re) : $signed(_GEN_5620); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5622 = 7'h30 == _T_9 ? $signed(regsB_82_re) : $signed(_GEN_5621); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5623 = 7'h31 == _T_9 ? $signed(regsB_92_re) : $signed(_GEN_5622); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5624 = 7'h32 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5623); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5625 = 7'h33 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5624); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5626 = 7'h34 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5625); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5627 = 7'h35 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5626); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5628 = 7'h36 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5627); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5629 = 7'h37 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5628); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5630 = 7'h38 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5629); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5631 = 7'h39 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5630); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5632 = 7'h3a == _T_9 ? $signed(32'sh0) : $signed(_GEN_5631); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5633 = 7'h3b == _T_9 ? $signed(32'sh0) : $signed(_GEN_5632); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5634 = 7'h3c == _T_9 ? $signed(regsB_3_re) : $signed(_GEN_5633); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5635 = 7'h3d == _T_9 ? $signed(regsB_13_re) : $signed(_GEN_5634); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5636 = 7'h3e == _T_9 ? $signed(regsB_23_re) : $signed(_GEN_5635); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5637 = 7'h3f == _T_9 ? $signed(regsB_33_re) : $signed(_GEN_5636); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5638 = 7'h40 == _T_9 ? $signed(regsB_43_re) : $signed(_GEN_5637); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5639 = 7'h41 == _T_9 ? $signed(regsB_53_re) : $signed(_GEN_5638); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5640 = 7'h42 == _T_9 ? $signed(regsB_63_re) : $signed(_GEN_5639); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5641 = 7'h43 == _T_9 ? $signed(regsB_73_re) : $signed(_GEN_5640); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5642 = 7'h44 == _T_9 ? $signed(regsB_83_re) : $signed(_GEN_5641); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5643 = 7'h45 == _T_9 ? $signed(regsB_93_re) : $signed(_GEN_5642); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5644 = 7'h46 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5643); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5645 = 7'h47 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5644); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5646 = 7'h48 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5645); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5647 = 7'h49 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5646); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5648 = 7'h4a == _T_9 ? $signed(32'sh0) : $signed(_GEN_5647); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5649 = 7'h4b == _T_9 ? $signed(32'sh0) : $signed(_GEN_5648); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5650 = 7'h4c == _T_9 ? $signed(32'sh0) : $signed(_GEN_5649); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5651 = 7'h4d == _T_9 ? $signed(32'sh0) : $signed(_GEN_5650); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5652 = 7'h4e == _T_9 ? $signed(32'sh0) : $signed(_GEN_5651); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5653 = 7'h4f == _T_9 ? $signed(32'sh0) : $signed(_GEN_5652); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5654 = 7'h50 == _T_9 ? $signed(regsB_4_re) : $signed(_GEN_5653); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5655 = 7'h51 == _T_9 ? $signed(regsB_14_re) : $signed(_GEN_5654); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5656 = 7'h52 == _T_9 ? $signed(regsB_24_re) : $signed(_GEN_5655); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5657 = 7'h53 == _T_9 ? $signed(regsB_34_re) : $signed(_GEN_5656); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5658 = 7'h54 == _T_9 ? $signed(regsB_44_re) : $signed(_GEN_5657); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5659 = 7'h55 == _T_9 ? $signed(regsB_54_re) : $signed(_GEN_5658); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5660 = 7'h56 == _T_9 ? $signed(regsB_64_re) : $signed(_GEN_5659); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5661 = 7'h57 == _T_9 ? $signed(regsB_74_re) : $signed(_GEN_5660); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5662 = 7'h58 == _T_9 ? $signed(regsB_84_re) : $signed(_GEN_5661); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5663 = 7'h59 == _T_9 ? $signed(regsB_94_re) : $signed(_GEN_5662); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5664 = 7'h5a == _T_9 ? $signed(32'sh0) : $signed(_GEN_5663); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5665 = 7'h5b == _T_9 ? $signed(32'sh0) : $signed(_GEN_5664); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5666 = 7'h5c == _T_9 ? $signed(32'sh0) : $signed(_GEN_5665); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5667 = 7'h5d == _T_9 ? $signed(32'sh0) : $signed(_GEN_5666); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5668 = 7'h5e == _T_9 ? $signed(32'sh0) : $signed(_GEN_5667); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5669 = 7'h5f == _T_9 ? $signed(32'sh0) : $signed(_GEN_5668); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5670 = 7'h60 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5669); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5671 = 7'h61 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5670); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5672 = 7'h62 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5671); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5673 = 7'h63 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5672); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5674 = 7'h64 == _T_9 ? $signed(regsB_5_re) : $signed(_GEN_5673); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5675 = 7'h65 == _T_9 ? $signed(regsB_15_re) : $signed(_GEN_5674); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5676 = 7'h66 == _T_9 ? $signed(regsB_25_re) : $signed(_GEN_5675); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5677 = 7'h67 == _T_9 ? $signed(regsB_35_re) : $signed(_GEN_5676); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5678 = 7'h68 == _T_9 ? $signed(regsB_45_re) : $signed(_GEN_5677); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5679 = 7'h69 == _T_9 ? $signed(regsB_55_re) : $signed(_GEN_5678); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5680 = 7'h6a == _T_9 ? $signed(regsB_65_re) : $signed(_GEN_5679); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5681 = 7'h6b == _T_9 ? $signed(regsB_75_re) : $signed(_GEN_5680); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5682 = 7'h6c == _T_9 ? $signed(regsB_85_re) : $signed(_GEN_5681); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5683 = 7'h6d == _T_9 ? $signed(regsB_95_re) : $signed(_GEN_5682); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5684 = 7'h6e == _T_9 ? $signed(32'sh0) : $signed(_GEN_5683); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5685 = 7'h6f == _T_9 ? $signed(32'sh0) : $signed(_GEN_5684); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5686 = 7'h70 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5685); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5687 = 7'h71 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5686); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5688 = 7'h72 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5687); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5689 = 7'h73 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5688); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5690 = 7'h74 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5689); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5691 = 7'h75 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5690); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5692 = 7'h76 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5691); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5693 = 7'h77 == _T_9 ? $signed(32'sh0) : $signed(_GEN_5692); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5694 = 7'h78 == _T_9 ? $signed(regsB_6_re) : $signed(_GEN_5693); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5695 = 7'h79 == _T_9 ? $signed(regsB_16_re) : $signed(_GEN_5694); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5696 = 7'h7a == _T_9 ? $signed(regsB_26_re) : $signed(_GEN_5695); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5697 = 7'h7b == _T_9 ? $signed(regsB_36_re) : $signed(_GEN_5696); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5698 = 7'h7c == _T_9 ? $signed(regsB_46_re) : $signed(_GEN_5697); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5699 = 7'h7d == _T_9 ? $signed(regsB_56_re) : $signed(_GEN_5698); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5700 = 7'h7e == _T_9 ? $signed(regsB_66_re) : $signed(_GEN_5699); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5701 = 7'h7f == _T_9 ? $signed(regsB_76_re) : $signed(_GEN_5700); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5702 = 8'h80 == _GEN_8950 ? $signed(regsB_86_re) : $signed(_GEN_5701); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5703 = 8'h81 == _GEN_8950 ? $signed(regsB_96_re) : $signed(_GEN_5702); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5704 = 8'h82 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5703); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5705 = 8'h83 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5704); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5706 = 8'h84 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5705); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5707 = 8'h85 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5706); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5708 = 8'h86 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5707); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5709 = 8'h87 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5708); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5710 = 8'h88 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5709); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5711 = 8'h89 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5710); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5712 = 8'h8a == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5711); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5713 = 8'h8b == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5712); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5714 = 8'h8c == _GEN_8950 ? $signed(regsB_7_re) : $signed(_GEN_5713); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5715 = 8'h8d == _GEN_8950 ? $signed(regsB_17_re) : $signed(_GEN_5714); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5716 = 8'h8e == _GEN_8950 ? $signed(regsB_27_re) : $signed(_GEN_5715); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5717 = 8'h8f == _GEN_8950 ? $signed(regsB_37_re) : $signed(_GEN_5716); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5718 = 8'h90 == _GEN_8950 ? $signed(regsB_47_re) : $signed(_GEN_5717); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5719 = 8'h91 == _GEN_8950 ? $signed(regsB_57_re) : $signed(_GEN_5718); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5720 = 8'h92 == _GEN_8950 ? $signed(regsB_67_re) : $signed(_GEN_5719); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5721 = 8'h93 == _GEN_8950 ? $signed(regsB_77_re) : $signed(_GEN_5720); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5722 = 8'h94 == _GEN_8950 ? $signed(regsB_87_re) : $signed(_GEN_5721); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5723 = 8'h95 == _GEN_8950 ? $signed(regsB_97_re) : $signed(_GEN_5722); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5724 = 8'h96 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5723); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5725 = 8'h97 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5724); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5726 = 8'h98 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5725); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5727 = 8'h99 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5726); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5728 = 8'h9a == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5727); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5729 = 8'h9b == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5728); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5730 = 8'h9c == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5729); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5731 = 8'h9d == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5730); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5732 = 8'h9e == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5731); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5733 = 8'h9f == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5732); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5734 = 8'ha0 == _GEN_8950 ? $signed(regsB_8_re) : $signed(_GEN_5733); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5735 = 8'ha1 == _GEN_8950 ? $signed(regsB_18_re) : $signed(_GEN_5734); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5736 = 8'ha2 == _GEN_8950 ? $signed(regsB_28_re) : $signed(_GEN_5735); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5737 = 8'ha3 == _GEN_8950 ? $signed(regsB_38_re) : $signed(_GEN_5736); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5738 = 8'ha4 == _GEN_8950 ? $signed(regsB_48_re) : $signed(_GEN_5737); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5739 = 8'ha5 == _GEN_8950 ? $signed(regsB_58_re) : $signed(_GEN_5738); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5740 = 8'ha6 == _GEN_8950 ? $signed(regsB_68_re) : $signed(_GEN_5739); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5741 = 8'ha7 == _GEN_8950 ? $signed(regsB_78_re) : $signed(_GEN_5740); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5742 = 8'ha8 == _GEN_8950 ? $signed(regsB_88_re) : $signed(_GEN_5741); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5743 = 8'ha9 == _GEN_8950 ? $signed(regsB_98_re) : $signed(_GEN_5742); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5744 = 8'haa == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5743); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5745 = 8'hab == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5744); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5746 = 8'hac == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5745); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5747 = 8'had == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5746); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5748 = 8'hae == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5747); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5749 = 8'haf == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5748); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5750 = 8'hb0 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5749); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5751 = 8'hb1 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5750); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5752 = 8'hb2 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5751); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5753 = 8'hb3 == _GEN_8950 ? $signed(32'sh0) : $signed(_GEN_5752); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5754 = 8'hb4 == _GEN_8950 ? $signed(regsB_9_re) : $signed(_GEN_5753); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5755 = 8'hb5 == _GEN_8950 ? $signed(regsB_19_re) : $signed(_GEN_5754); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5756 = 8'hb6 == _GEN_8950 ? $signed(regsB_29_re) : $signed(_GEN_5755); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5757 = 8'hb7 == _GEN_8950 ? $signed(regsB_39_re) : $signed(_GEN_5756); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5758 = 8'hb8 == _GEN_8950 ? $signed(regsB_49_re) : $signed(_GEN_5757); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5759 = 8'hb9 == _GEN_8950 ? $signed(regsB_59_re) : $signed(_GEN_5758); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5760 = 8'hba == _GEN_8950 ? $signed(regsB_69_re) : $signed(_GEN_5759); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5761 = 8'hbb == _GEN_8950 ? $signed(regsB_79_re) : $signed(_GEN_5760); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5762 = 8'hbc == _GEN_8950 ? $signed(regsB_89_re) : $signed(_GEN_5761); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5763 = 8'hbd == _GEN_8950 ? $signed(regsB_99_re) : $signed(_GEN_5762); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5765 = 7'h1 == _T_12 ? $signed(regsB_10_im) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5766 = 7'h2 == _T_12 ? $signed(regsB_20_im) : $signed(_GEN_5765); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5767 = 7'h3 == _T_12 ? $signed(regsB_30_im) : $signed(_GEN_5766); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5768 = 7'h4 == _T_12 ? $signed(regsB_40_im) : $signed(_GEN_5767); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5769 = 7'h5 == _T_12 ? $signed(regsB_50_im) : $signed(_GEN_5768); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5770 = 7'h6 == _T_12 ? $signed(regsB_60_im) : $signed(_GEN_5769); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5771 = 7'h7 == _T_12 ? $signed(regsB_70_im) : $signed(_GEN_5770); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5772 = 7'h8 == _T_12 ? $signed(regsB_80_im) : $signed(_GEN_5771); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5773 = 7'h9 == _T_12 ? $signed(regsB_90_im) : $signed(_GEN_5772); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5774 = 7'ha == _T_12 ? $signed(32'sh0) : $signed(_GEN_5773); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5775 = 7'hb == _T_12 ? $signed(32'sh0) : $signed(_GEN_5774); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5776 = 7'hc == _T_12 ? $signed(32'sh0) : $signed(_GEN_5775); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5777 = 7'hd == _T_12 ? $signed(32'sh0) : $signed(_GEN_5776); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5778 = 7'he == _T_12 ? $signed(32'sh0) : $signed(_GEN_5777); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5779 = 7'hf == _T_12 ? $signed(32'sh0) : $signed(_GEN_5778); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5780 = 7'h10 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5779); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5781 = 7'h11 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5780); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5782 = 7'h12 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5781); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5783 = 7'h13 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5782); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5784 = 7'h14 == _T_12 ? $signed(regsB_1_im) : $signed(_GEN_5783); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5785 = 7'h15 == _T_12 ? $signed(regsB_11_im) : $signed(_GEN_5784); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5786 = 7'h16 == _T_12 ? $signed(regsB_21_im) : $signed(_GEN_5785); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5787 = 7'h17 == _T_12 ? $signed(regsB_31_im) : $signed(_GEN_5786); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5788 = 7'h18 == _T_12 ? $signed(regsB_41_im) : $signed(_GEN_5787); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5789 = 7'h19 == _T_12 ? $signed(regsB_51_im) : $signed(_GEN_5788); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5790 = 7'h1a == _T_12 ? $signed(regsB_61_im) : $signed(_GEN_5789); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5791 = 7'h1b == _T_12 ? $signed(regsB_71_im) : $signed(_GEN_5790); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5792 = 7'h1c == _T_12 ? $signed(regsB_81_im) : $signed(_GEN_5791); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5793 = 7'h1d == _T_12 ? $signed(regsB_91_im) : $signed(_GEN_5792); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5794 = 7'h1e == _T_12 ? $signed(32'sh0) : $signed(_GEN_5793); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5795 = 7'h1f == _T_12 ? $signed(32'sh0) : $signed(_GEN_5794); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5796 = 7'h20 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5795); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5797 = 7'h21 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5796); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5798 = 7'h22 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5797); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5799 = 7'h23 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5798); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5800 = 7'h24 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5799); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5801 = 7'h25 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5800); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5802 = 7'h26 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5801); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5803 = 7'h27 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5802); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5804 = 7'h28 == _T_12 ? $signed(regsB_2_im) : $signed(_GEN_5803); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5805 = 7'h29 == _T_12 ? $signed(regsB_12_im) : $signed(_GEN_5804); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5806 = 7'h2a == _T_12 ? $signed(regsB_22_im) : $signed(_GEN_5805); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5807 = 7'h2b == _T_12 ? $signed(regsB_32_im) : $signed(_GEN_5806); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5808 = 7'h2c == _T_12 ? $signed(regsB_42_im) : $signed(_GEN_5807); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5809 = 7'h2d == _T_12 ? $signed(regsB_52_im) : $signed(_GEN_5808); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5810 = 7'h2e == _T_12 ? $signed(regsB_62_im) : $signed(_GEN_5809); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5811 = 7'h2f == _T_12 ? $signed(regsB_72_im) : $signed(_GEN_5810); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5812 = 7'h30 == _T_12 ? $signed(regsB_82_im) : $signed(_GEN_5811); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5813 = 7'h31 == _T_12 ? $signed(regsB_92_im) : $signed(_GEN_5812); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5814 = 7'h32 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5813); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5815 = 7'h33 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5814); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5816 = 7'h34 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5815); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5817 = 7'h35 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5816); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5818 = 7'h36 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5817); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5819 = 7'h37 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5818); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5820 = 7'h38 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5819); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5821 = 7'h39 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5820); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5822 = 7'h3a == _T_12 ? $signed(32'sh0) : $signed(_GEN_5821); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5823 = 7'h3b == _T_12 ? $signed(32'sh0) : $signed(_GEN_5822); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5824 = 7'h3c == _T_12 ? $signed(regsB_3_im) : $signed(_GEN_5823); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5825 = 7'h3d == _T_12 ? $signed(regsB_13_im) : $signed(_GEN_5824); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5826 = 7'h3e == _T_12 ? $signed(regsB_23_im) : $signed(_GEN_5825); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5827 = 7'h3f == _T_12 ? $signed(regsB_33_im) : $signed(_GEN_5826); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5828 = 7'h40 == _T_12 ? $signed(regsB_43_im) : $signed(_GEN_5827); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5829 = 7'h41 == _T_12 ? $signed(regsB_53_im) : $signed(_GEN_5828); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5830 = 7'h42 == _T_12 ? $signed(regsB_63_im) : $signed(_GEN_5829); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5831 = 7'h43 == _T_12 ? $signed(regsB_73_im) : $signed(_GEN_5830); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5832 = 7'h44 == _T_12 ? $signed(regsB_83_im) : $signed(_GEN_5831); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5833 = 7'h45 == _T_12 ? $signed(regsB_93_im) : $signed(_GEN_5832); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5834 = 7'h46 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5833); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5835 = 7'h47 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5834); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5836 = 7'h48 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5835); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5837 = 7'h49 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5836); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5838 = 7'h4a == _T_12 ? $signed(32'sh0) : $signed(_GEN_5837); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5839 = 7'h4b == _T_12 ? $signed(32'sh0) : $signed(_GEN_5838); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5840 = 7'h4c == _T_12 ? $signed(32'sh0) : $signed(_GEN_5839); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5841 = 7'h4d == _T_12 ? $signed(32'sh0) : $signed(_GEN_5840); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5842 = 7'h4e == _T_12 ? $signed(32'sh0) : $signed(_GEN_5841); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5843 = 7'h4f == _T_12 ? $signed(32'sh0) : $signed(_GEN_5842); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5844 = 7'h50 == _T_12 ? $signed(regsB_4_im) : $signed(_GEN_5843); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5845 = 7'h51 == _T_12 ? $signed(regsB_14_im) : $signed(_GEN_5844); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5846 = 7'h52 == _T_12 ? $signed(regsB_24_im) : $signed(_GEN_5845); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5847 = 7'h53 == _T_12 ? $signed(regsB_34_im) : $signed(_GEN_5846); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5848 = 7'h54 == _T_12 ? $signed(regsB_44_im) : $signed(_GEN_5847); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5849 = 7'h55 == _T_12 ? $signed(regsB_54_im) : $signed(_GEN_5848); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5850 = 7'h56 == _T_12 ? $signed(regsB_64_im) : $signed(_GEN_5849); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5851 = 7'h57 == _T_12 ? $signed(regsB_74_im) : $signed(_GEN_5850); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5852 = 7'h58 == _T_12 ? $signed(regsB_84_im) : $signed(_GEN_5851); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5853 = 7'h59 == _T_12 ? $signed(regsB_94_im) : $signed(_GEN_5852); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5854 = 7'h5a == _T_12 ? $signed(32'sh0) : $signed(_GEN_5853); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5855 = 7'h5b == _T_12 ? $signed(32'sh0) : $signed(_GEN_5854); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5856 = 7'h5c == _T_12 ? $signed(32'sh0) : $signed(_GEN_5855); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5857 = 7'h5d == _T_12 ? $signed(32'sh0) : $signed(_GEN_5856); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5858 = 7'h5e == _T_12 ? $signed(32'sh0) : $signed(_GEN_5857); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5859 = 7'h5f == _T_12 ? $signed(32'sh0) : $signed(_GEN_5858); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5860 = 7'h60 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5859); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5861 = 7'h61 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5860); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5862 = 7'h62 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5861); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5863 = 7'h63 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5862); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5864 = 7'h64 == _T_12 ? $signed(regsB_5_im) : $signed(_GEN_5863); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5865 = 7'h65 == _T_12 ? $signed(regsB_15_im) : $signed(_GEN_5864); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5866 = 7'h66 == _T_12 ? $signed(regsB_25_im) : $signed(_GEN_5865); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5867 = 7'h67 == _T_12 ? $signed(regsB_35_im) : $signed(_GEN_5866); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5868 = 7'h68 == _T_12 ? $signed(regsB_45_im) : $signed(_GEN_5867); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5869 = 7'h69 == _T_12 ? $signed(regsB_55_im) : $signed(_GEN_5868); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5870 = 7'h6a == _T_12 ? $signed(regsB_65_im) : $signed(_GEN_5869); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5871 = 7'h6b == _T_12 ? $signed(regsB_75_im) : $signed(_GEN_5870); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5872 = 7'h6c == _T_12 ? $signed(regsB_85_im) : $signed(_GEN_5871); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5873 = 7'h6d == _T_12 ? $signed(regsB_95_im) : $signed(_GEN_5872); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5874 = 7'h6e == _T_12 ? $signed(32'sh0) : $signed(_GEN_5873); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5875 = 7'h6f == _T_12 ? $signed(32'sh0) : $signed(_GEN_5874); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5876 = 7'h70 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5875); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5877 = 7'h71 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5876); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5878 = 7'h72 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5877); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5879 = 7'h73 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5878); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5880 = 7'h74 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5879); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5881 = 7'h75 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5880); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5882 = 7'h76 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5881); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5883 = 7'h77 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5882); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5884 = 7'h78 == _T_12 ? $signed(regsB_6_im) : $signed(_GEN_5883); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5885 = 7'h79 == _T_12 ? $signed(regsB_16_im) : $signed(_GEN_5884); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5886 = 7'h7a == _T_12 ? $signed(regsB_26_im) : $signed(_GEN_5885); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5887 = 7'h7b == _T_12 ? $signed(regsB_36_im) : $signed(_GEN_5886); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5888 = 7'h7c == _T_12 ? $signed(regsB_46_im) : $signed(_GEN_5887); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5889 = 7'h7d == _T_12 ? $signed(regsB_56_im) : $signed(_GEN_5888); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5890 = 7'h7e == _T_12 ? $signed(regsB_66_im) : $signed(_GEN_5889); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5891 = 7'h7f == _T_12 ? $signed(regsB_76_im) : $signed(_GEN_5890); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5892 = 8'h80 == _GEN_9075 ? $signed(regsB_86_im) : $signed(_GEN_5891); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5893 = 8'h81 == _GEN_9075 ? $signed(regsB_96_im) : $signed(_GEN_5892); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5894 = 8'h82 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5893); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5895 = 8'h83 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5894); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5896 = 8'h84 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5895); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5897 = 8'h85 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5896); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5898 = 8'h86 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5897); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5899 = 8'h87 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5898); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5900 = 8'h88 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5899); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5901 = 8'h89 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5900); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5902 = 8'h8a == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5901); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5903 = 8'h8b == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5902); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5904 = 8'h8c == _GEN_9075 ? $signed(regsB_7_im) : $signed(_GEN_5903); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5905 = 8'h8d == _GEN_9075 ? $signed(regsB_17_im) : $signed(_GEN_5904); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5906 = 8'h8e == _GEN_9075 ? $signed(regsB_27_im) : $signed(_GEN_5905); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5907 = 8'h8f == _GEN_9075 ? $signed(regsB_37_im) : $signed(_GEN_5906); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5908 = 8'h90 == _GEN_9075 ? $signed(regsB_47_im) : $signed(_GEN_5907); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5909 = 8'h91 == _GEN_9075 ? $signed(regsB_57_im) : $signed(_GEN_5908); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5910 = 8'h92 == _GEN_9075 ? $signed(regsB_67_im) : $signed(_GEN_5909); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5911 = 8'h93 == _GEN_9075 ? $signed(regsB_77_im) : $signed(_GEN_5910); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5912 = 8'h94 == _GEN_9075 ? $signed(regsB_87_im) : $signed(_GEN_5911); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5913 = 8'h95 == _GEN_9075 ? $signed(regsB_97_im) : $signed(_GEN_5912); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5914 = 8'h96 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5913); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5915 = 8'h97 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5914); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5916 = 8'h98 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5915); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5917 = 8'h99 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5916); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5918 = 8'h9a == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5917); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5919 = 8'h9b == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5918); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5920 = 8'h9c == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5919); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5921 = 8'h9d == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5920); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5922 = 8'h9e == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5921); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5923 = 8'h9f == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5922); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5924 = 8'ha0 == _GEN_9075 ? $signed(regsB_8_im) : $signed(_GEN_5923); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5925 = 8'ha1 == _GEN_9075 ? $signed(regsB_18_im) : $signed(_GEN_5924); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5926 = 8'ha2 == _GEN_9075 ? $signed(regsB_28_im) : $signed(_GEN_5925); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5927 = 8'ha3 == _GEN_9075 ? $signed(regsB_38_im) : $signed(_GEN_5926); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5928 = 8'ha4 == _GEN_9075 ? $signed(regsB_48_im) : $signed(_GEN_5927); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5929 = 8'ha5 == _GEN_9075 ? $signed(regsB_58_im) : $signed(_GEN_5928); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5930 = 8'ha6 == _GEN_9075 ? $signed(regsB_68_im) : $signed(_GEN_5929); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5931 = 8'ha7 == _GEN_9075 ? $signed(regsB_78_im) : $signed(_GEN_5930); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5932 = 8'ha8 == _GEN_9075 ? $signed(regsB_88_im) : $signed(_GEN_5931); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5933 = 8'ha9 == _GEN_9075 ? $signed(regsB_98_im) : $signed(_GEN_5932); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5934 = 8'haa == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5933); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5935 = 8'hab == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5934); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5936 = 8'hac == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5935); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5937 = 8'had == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5936); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5938 = 8'hae == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5937); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5939 = 8'haf == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5938); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5940 = 8'hb0 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5939); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5941 = 8'hb1 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5940); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5942 = 8'hb2 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5941); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5943 = 8'hb3 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_5942); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5944 = 8'hb4 == _GEN_9075 ? $signed(regsB_9_im) : $signed(_GEN_5943); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5945 = 8'hb5 == _GEN_9075 ? $signed(regsB_19_im) : $signed(_GEN_5944); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5946 = 8'hb6 == _GEN_9075 ? $signed(regsB_29_im) : $signed(_GEN_5945); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5947 = 8'hb7 == _GEN_9075 ? $signed(regsB_39_im) : $signed(_GEN_5946); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5948 = 8'hb8 == _GEN_9075 ? $signed(regsB_49_im) : $signed(_GEN_5947); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5949 = 8'hb9 == _GEN_9075 ? $signed(regsB_59_im) : $signed(_GEN_5948); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5950 = 8'hba == _GEN_9075 ? $signed(regsB_69_im) : $signed(_GEN_5949); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5951 = 8'hbb == _GEN_9075 ? $signed(regsB_79_im) : $signed(_GEN_5950); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5952 = 8'hbc == _GEN_9075 ? $signed(regsB_89_im) : $signed(_GEN_5951); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5953 = 8'hbd == _GEN_9075 ? $signed(regsB_99_im) : $signed(_GEN_5952); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5955 = 7'h1 == _T_12 ? $signed(regsB_10_re) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5956 = 7'h2 == _T_12 ? $signed(regsB_20_re) : $signed(_GEN_5955); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5957 = 7'h3 == _T_12 ? $signed(regsB_30_re) : $signed(_GEN_5956); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5958 = 7'h4 == _T_12 ? $signed(regsB_40_re) : $signed(_GEN_5957); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5959 = 7'h5 == _T_12 ? $signed(regsB_50_re) : $signed(_GEN_5958); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5960 = 7'h6 == _T_12 ? $signed(regsB_60_re) : $signed(_GEN_5959); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5961 = 7'h7 == _T_12 ? $signed(regsB_70_re) : $signed(_GEN_5960); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5962 = 7'h8 == _T_12 ? $signed(regsB_80_re) : $signed(_GEN_5961); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5963 = 7'h9 == _T_12 ? $signed(regsB_90_re) : $signed(_GEN_5962); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5964 = 7'ha == _T_12 ? $signed(32'sh0) : $signed(_GEN_5963); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5965 = 7'hb == _T_12 ? $signed(32'sh0) : $signed(_GEN_5964); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5966 = 7'hc == _T_12 ? $signed(32'sh0) : $signed(_GEN_5965); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5967 = 7'hd == _T_12 ? $signed(32'sh0) : $signed(_GEN_5966); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5968 = 7'he == _T_12 ? $signed(32'sh0) : $signed(_GEN_5967); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5969 = 7'hf == _T_12 ? $signed(32'sh0) : $signed(_GEN_5968); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5970 = 7'h10 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5969); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5971 = 7'h11 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5970); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5972 = 7'h12 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5971); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5973 = 7'h13 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5972); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5974 = 7'h14 == _T_12 ? $signed(regsB_1_re) : $signed(_GEN_5973); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5975 = 7'h15 == _T_12 ? $signed(regsB_11_re) : $signed(_GEN_5974); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5976 = 7'h16 == _T_12 ? $signed(regsB_21_re) : $signed(_GEN_5975); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5977 = 7'h17 == _T_12 ? $signed(regsB_31_re) : $signed(_GEN_5976); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5978 = 7'h18 == _T_12 ? $signed(regsB_41_re) : $signed(_GEN_5977); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5979 = 7'h19 == _T_12 ? $signed(regsB_51_re) : $signed(_GEN_5978); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5980 = 7'h1a == _T_12 ? $signed(regsB_61_re) : $signed(_GEN_5979); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5981 = 7'h1b == _T_12 ? $signed(regsB_71_re) : $signed(_GEN_5980); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5982 = 7'h1c == _T_12 ? $signed(regsB_81_re) : $signed(_GEN_5981); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5983 = 7'h1d == _T_12 ? $signed(regsB_91_re) : $signed(_GEN_5982); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5984 = 7'h1e == _T_12 ? $signed(32'sh0) : $signed(_GEN_5983); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5985 = 7'h1f == _T_12 ? $signed(32'sh0) : $signed(_GEN_5984); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5986 = 7'h20 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5985); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5987 = 7'h21 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5986); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5988 = 7'h22 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5987); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5989 = 7'h23 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5988); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5990 = 7'h24 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5989); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5991 = 7'h25 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5990); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5992 = 7'h26 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5991); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5993 = 7'h27 == _T_12 ? $signed(32'sh0) : $signed(_GEN_5992); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5994 = 7'h28 == _T_12 ? $signed(regsB_2_re) : $signed(_GEN_5993); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5995 = 7'h29 == _T_12 ? $signed(regsB_12_re) : $signed(_GEN_5994); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5996 = 7'h2a == _T_12 ? $signed(regsB_22_re) : $signed(_GEN_5995); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5997 = 7'h2b == _T_12 ? $signed(regsB_32_re) : $signed(_GEN_5996); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5998 = 7'h2c == _T_12 ? $signed(regsB_42_re) : $signed(_GEN_5997); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_5999 = 7'h2d == _T_12 ? $signed(regsB_52_re) : $signed(_GEN_5998); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6000 = 7'h2e == _T_12 ? $signed(regsB_62_re) : $signed(_GEN_5999); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6001 = 7'h2f == _T_12 ? $signed(regsB_72_re) : $signed(_GEN_6000); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6002 = 7'h30 == _T_12 ? $signed(regsB_82_re) : $signed(_GEN_6001); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6003 = 7'h31 == _T_12 ? $signed(regsB_92_re) : $signed(_GEN_6002); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6004 = 7'h32 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6003); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6005 = 7'h33 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6004); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6006 = 7'h34 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6005); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6007 = 7'h35 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6006); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6008 = 7'h36 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6007); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6009 = 7'h37 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6008); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6010 = 7'h38 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6009); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6011 = 7'h39 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6010); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6012 = 7'h3a == _T_12 ? $signed(32'sh0) : $signed(_GEN_6011); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6013 = 7'h3b == _T_12 ? $signed(32'sh0) : $signed(_GEN_6012); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6014 = 7'h3c == _T_12 ? $signed(regsB_3_re) : $signed(_GEN_6013); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6015 = 7'h3d == _T_12 ? $signed(regsB_13_re) : $signed(_GEN_6014); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6016 = 7'h3e == _T_12 ? $signed(regsB_23_re) : $signed(_GEN_6015); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6017 = 7'h3f == _T_12 ? $signed(regsB_33_re) : $signed(_GEN_6016); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6018 = 7'h40 == _T_12 ? $signed(regsB_43_re) : $signed(_GEN_6017); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6019 = 7'h41 == _T_12 ? $signed(regsB_53_re) : $signed(_GEN_6018); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6020 = 7'h42 == _T_12 ? $signed(regsB_63_re) : $signed(_GEN_6019); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6021 = 7'h43 == _T_12 ? $signed(regsB_73_re) : $signed(_GEN_6020); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6022 = 7'h44 == _T_12 ? $signed(regsB_83_re) : $signed(_GEN_6021); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6023 = 7'h45 == _T_12 ? $signed(regsB_93_re) : $signed(_GEN_6022); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6024 = 7'h46 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6023); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6025 = 7'h47 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6024); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6026 = 7'h48 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6025); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6027 = 7'h49 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6026); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6028 = 7'h4a == _T_12 ? $signed(32'sh0) : $signed(_GEN_6027); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6029 = 7'h4b == _T_12 ? $signed(32'sh0) : $signed(_GEN_6028); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6030 = 7'h4c == _T_12 ? $signed(32'sh0) : $signed(_GEN_6029); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6031 = 7'h4d == _T_12 ? $signed(32'sh0) : $signed(_GEN_6030); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6032 = 7'h4e == _T_12 ? $signed(32'sh0) : $signed(_GEN_6031); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6033 = 7'h4f == _T_12 ? $signed(32'sh0) : $signed(_GEN_6032); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6034 = 7'h50 == _T_12 ? $signed(regsB_4_re) : $signed(_GEN_6033); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6035 = 7'h51 == _T_12 ? $signed(regsB_14_re) : $signed(_GEN_6034); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6036 = 7'h52 == _T_12 ? $signed(regsB_24_re) : $signed(_GEN_6035); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6037 = 7'h53 == _T_12 ? $signed(regsB_34_re) : $signed(_GEN_6036); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6038 = 7'h54 == _T_12 ? $signed(regsB_44_re) : $signed(_GEN_6037); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6039 = 7'h55 == _T_12 ? $signed(regsB_54_re) : $signed(_GEN_6038); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6040 = 7'h56 == _T_12 ? $signed(regsB_64_re) : $signed(_GEN_6039); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6041 = 7'h57 == _T_12 ? $signed(regsB_74_re) : $signed(_GEN_6040); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6042 = 7'h58 == _T_12 ? $signed(regsB_84_re) : $signed(_GEN_6041); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6043 = 7'h59 == _T_12 ? $signed(regsB_94_re) : $signed(_GEN_6042); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6044 = 7'h5a == _T_12 ? $signed(32'sh0) : $signed(_GEN_6043); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6045 = 7'h5b == _T_12 ? $signed(32'sh0) : $signed(_GEN_6044); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6046 = 7'h5c == _T_12 ? $signed(32'sh0) : $signed(_GEN_6045); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6047 = 7'h5d == _T_12 ? $signed(32'sh0) : $signed(_GEN_6046); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6048 = 7'h5e == _T_12 ? $signed(32'sh0) : $signed(_GEN_6047); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6049 = 7'h5f == _T_12 ? $signed(32'sh0) : $signed(_GEN_6048); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6050 = 7'h60 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6049); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6051 = 7'h61 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6050); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6052 = 7'h62 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6051); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6053 = 7'h63 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6052); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6054 = 7'h64 == _T_12 ? $signed(regsB_5_re) : $signed(_GEN_6053); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6055 = 7'h65 == _T_12 ? $signed(regsB_15_re) : $signed(_GEN_6054); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6056 = 7'h66 == _T_12 ? $signed(regsB_25_re) : $signed(_GEN_6055); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6057 = 7'h67 == _T_12 ? $signed(regsB_35_re) : $signed(_GEN_6056); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6058 = 7'h68 == _T_12 ? $signed(regsB_45_re) : $signed(_GEN_6057); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6059 = 7'h69 == _T_12 ? $signed(regsB_55_re) : $signed(_GEN_6058); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6060 = 7'h6a == _T_12 ? $signed(regsB_65_re) : $signed(_GEN_6059); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6061 = 7'h6b == _T_12 ? $signed(regsB_75_re) : $signed(_GEN_6060); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6062 = 7'h6c == _T_12 ? $signed(regsB_85_re) : $signed(_GEN_6061); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6063 = 7'h6d == _T_12 ? $signed(regsB_95_re) : $signed(_GEN_6062); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6064 = 7'h6e == _T_12 ? $signed(32'sh0) : $signed(_GEN_6063); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6065 = 7'h6f == _T_12 ? $signed(32'sh0) : $signed(_GEN_6064); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6066 = 7'h70 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6065); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6067 = 7'h71 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6066); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6068 = 7'h72 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6067); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6069 = 7'h73 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6068); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6070 = 7'h74 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6069); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6071 = 7'h75 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6070); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6072 = 7'h76 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6071); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6073 = 7'h77 == _T_12 ? $signed(32'sh0) : $signed(_GEN_6072); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6074 = 7'h78 == _T_12 ? $signed(regsB_6_re) : $signed(_GEN_6073); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6075 = 7'h79 == _T_12 ? $signed(regsB_16_re) : $signed(_GEN_6074); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6076 = 7'h7a == _T_12 ? $signed(regsB_26_re) : $signed(_GEN_6075); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6077 = 7'h7b == _T_12 ? $signed(regsB_36_re) : $signed(_GEN_6076); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6078 = 7'h7c == _T_12 ? $signed(regsB_46_re) : $signed(_GEN_6077); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6079 = 7'h7d == _T_12 ? $signed(regsB_56_re) : $signed(_GEN_6078); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6080 = 7'h7e == _T_12 ? $signed(regsB_66_re) : $signed(_GEN_6079); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6081 = 7'h7f == _T_12 ? $signed(regsB_76_re) : $signed(_GEN_6080); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6082 = 8'h80 == _GEN_9075 ? $signed(regsB_86_re) : $signed(_GEN_6081); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6083 = 8'h81 == _GEN_9075 ? $signed(regsB_96_re) : $signed(_GEN_6082); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6084 = 8'h82 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6083); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6085 = 8'h83 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6084); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6086 = 8'h84 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6085); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6087 = 8'h85 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6086); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6088 = 8'h86 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6087); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6089 = 8'h87 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6088); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6090 = 8'h88 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6089); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6091 = 8'h89 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6090); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6092 = 8'h8a == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6091); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6093 = 8'h8b == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6092); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6094 = 8'h8c == _GEN_9075 ? $signed(regsB_7_re) : $signed(_GEN_6093); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6095 = 8'h8d == _GEN_9075 ? $signed(regsB_17_re) : $signed(_GEN_6094); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6096 = 8'h8e == _GEN_9075 ? $signed(regsB_27_re) : $signed(_GEN_6095); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6097 = 8'h8f == _GEN_9075 ? $signed(regsB_37_re) : $signed(_GEN_6096); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6098 = 8'h90 == _GEN_9075 ? $signed(regsB_47_re) : $signed(_GEN_6097); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6099 = 8'h91 == _GEN_9075 ? $signed(regsB_57_re) : $signed(_GEN_6098); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6100 = 8'h92 == _GEN_9075 ? $signed(regsB_67_re) : $signed(_GEN_6099); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6101 = 8'h93 == _GEN_9075 ? $signed(regsB_77_re) : $signed(_GEN_6100); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6102 = 8'h94 == _GEN_9075 ? $signed(regsB_87_re) : $signed(_GEN_6101); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6103 = 8'h95 == _GEN_9075 ? $signed(regsB_97_re) : $signed(_GEN_6102); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6104 = 8'h96 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6103); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6105 = 8'h97 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6104); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6106 = 8'h98 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6105); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6107 = 8'h99 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6106); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6108 = 8'h9a == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6107); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6109 = 8'h9b == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6108); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6110 = 8'h9c == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6109); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6111 = 8'h9d == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6110); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6112 = 8'h9e == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6111); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6113 = 8'h9f == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6112); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6114 = 8'ha0 == _GEN_9075 ? $signed(regsB_8_re) : $signed(_GEN_6113); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6115 = 8'ha1 == _GEN_9075 ? $signed(regsB_18_re) : $signed(_GEN_6114); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6116 = 8'ha2 == _GEN_9075 ? $signed(regsB_28_re) : $signed(_GEN_6115); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6117 = 8'ha3 == _GEN_9075 ? $signed(regsB_38_re) : $signed(_GEN_6116); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6118 = 8'ha4 == _GEN_9075 ? $signed(regsB_48_re) : $signed(_GEN_6117); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6119 = 8'ha5 == _GEN_9075 ? $signed(regsB_58_re) : $signed(_GEN_6118); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6120 = 8'ha6 == _GEN_9075 ? $signed(regsB_68_re) : $signed(_GEN_6119); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6121 = 8'ha7 == _GEN_9075 ? $signed(regsB_78_re) : $signed(_GEN_6120); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6122 = 8'ha8 == _GEN_9075 ? $signed(regsB_88_re) : $signed(_GEN_6121); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6123 = 8'ha9 == _GEN_9075 ? $signed(regsB_98_re) : $signed(_GEN_6122); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6124 = 8'haa == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6123); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6125 = 8'hab == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6124); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6126 = 8'hac == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6125); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6127 = 8'had == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6126); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6128 = 8'hae == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6127); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6129 = 8'haf == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6128); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6130 = 8'hb0 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6129); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6131 = 8'hb1 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6130); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6132 = 8'hb2 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6131); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6133 = 8'hb3 == _GEN_9075 ? $signed(32'sh0) : $signed(_GEN_6132); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6134 = 8'hb4 == _GEN_9075 ? $signed(regsB_9_re) : $signed(_GEN_6133); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6135 = 8'hb5 == _GEN_9075 ? $signed(regsB_19_re) : $signed(_GEN_6134); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6136 = 8'hb6 == _GEN_9075 ? $signed(regsB_29_re) : $signed(_GEN_6135); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6137 = 8'hb7 == _GEN_9075 ? $signed(regsB_39_re) : $signed(_GEN_6136); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6138 = 8'hb8 == _GEN_9075 ? $signed(regsB_49_re) : $signed(_GEN_6137); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6139 = 8'hb9 == _GEN_9075 ? $signed(regsB_59_re) : $signed(_GEN_6138); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6140 = 8'hba == _GEN_9075 ? $signed(regsB_69_re) : $signed(_GEN_6139); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6141 = 8'hbb == _GEN_9075 ? $signed(regsB_79_re) : $signed(_GEN_6140); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6142 = 8'hbc == _GEN_9075 ? $signed(regsB_89_re) : $signed(_GEN_6141); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6143 = 8'hbd == _GEN_9075 ? $signed(regsB_99_re) : $signed(_GEN_6142); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6145 = 8'h1 == _T_15 ? $signed(regsB_10_im) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6146 = 8'h2 == _T_15 ? $signed(regsB_20_im) : $signed(_GEN_6145); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6147 = 8'h3 == _T_15 ? $signed(regsB_30_im) : $signed(_GEN_6146); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6148 = 8'h4 == _T_15 ? $signed(regsB_40_im) : $signed(_GEN_6147); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6149 = 8'h5 == _T_15 ? $signed(regsB_50_im) : $signed(_GEN_6148); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6150 = 8'h6 == _T_15 ? $signed(regsB_60_im) : $signed(_GEN_6149); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6151 = 8'h7 == _T_15 ? $signed(regsB_70_im) : $signed(_GEN_6150); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6152 = 8'h8 == _T_15 ? $signed(regsB_80_im) : $signed(_GEN_6151); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6153 = 8'h9 == _T_15 ? $signed(regsB_90_im) : $signed(_GEN_6152); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6154 = 8'ha == _T_15 ? $signed(32'sh0) : $signed(_GEN_6153); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6155 = 8'hb == _T_15 ? $signed(32'sh0) : $signed(_GEN_6154); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6156 = 8'hc == _T_15 ? $signed(32'sh0) : $signed(_GEN_6155); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6157 = 8'hd == _T_15 ? $signed(32'sh0) : $signed(_GEN_6156); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6158 = 8'he == _T_15 ? $signed(32'sh0) : $signed(_GEN_6157); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6159 = 8'hf == _T_15 ? $signed(32'sh0) : $signed(_GEN_6158); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6160 = 8'h10 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6159); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6161 = 8'h11 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6160); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6162 = 8'h12 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6161); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6163 = 8'h13 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6162); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6164 = 8'h14 == _T_15 ? $signed(regsB_1_im) : $signed(_GEN_6163); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6165 = 8'h15 == _T_15 ? $signed(regsB_11_im) : $signed(_GEN_6164); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6166 = 8'h16 == _T_15 ? $signed(regsB_21_im) : $signed(_GEN_6165); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6167 = 8'h17 == _T_15 ? $signed(regsB_31_im) : $signed(_GEN_6166); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6168 = 8'h18 == _T_15 ? $signed(regsB_41_im) : $signed(_GEN_6167); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6169 = 8'h19 == _T_15 ? $signed(regsB_51_im) : $signed(_GEN_6168); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6170 = 8'h1a == _T_15 ? $signed(regsB_61_im) : $signed(_GEN_6169); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6171 = 8'h1b == _T_15 ? $signed(regsB_71_im) : $signed(_GEN_6170); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6172 = 8'h1c == _T_15 ? $signed(regsB_81_im) : $signed(_GEN_6171); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6173 = 8'h1d == _T_15 ? $signed(regsB_91_im) : $signed(_GEN_6172); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6174 = 8'h1e == _T_15 ? $signed(32'sh0) : $signed(_GEN_6173); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6175 = 8'h1f == _T_15 ? $signed(32'sh0) : $signed(_GEN_6174); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6176 = 8'h20 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6175); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6177 = 8'h21 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6176); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6178 = 8'h22 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6177); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6179 = 8'h23 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6178); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6180 = 8'h24 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6179); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6181 = 8'h25 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6180); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6182 = 8'h26 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6181); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6183 = 8'h27 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6182); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6184 = 8'h28 == _T_15 ? $signed(regsB_2_im) : $signed(_GEN_6183); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6185 = 8'h29 == _T_15 ? $signed(regsB_12_im) : $signed(_GEN_6184); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6186 = 8'h2a == _T_15 ? $signed(regsB_22_im) : $signed(_GEN_6185); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6187 = 8'h2b == _T_15 ? $signed(regsB_32_im) : $signed(_GEN_6186); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6188 = 8'h2c == _T_15 ? $signed(regsB_42_im) : $signed(_GEN_6187); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6189 = 8'h2d == _T_15 ? $signed(regsB_52_im) : $signed(_GEN_6188); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6190 = 8'h2e == _T_15 ? $signed(regsB_62_im) : $signed(_GEN_6189); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6191 = 8'h2f == _T_15 ? $signed(regsB_72_im) : $signed(_GEN_6190); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6192 = 8'h30 == _T_15 ? $signed(regsB_82_im) : $signed(_GEN_6191); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6193 = 8'h31 == _T_15 ? $signed(regsB_92_im) : $signed(_GEN_6192); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6194 = 8'h32 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6193); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6195 = 8'h33 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6194); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6196 = 8'h34 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6195); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6197 = 8'h35 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6196); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6198 = 8'h36 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6197); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6199 = 8'h37 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6198); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6200 = 8'h38 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6199); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6201 = 8'h39 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6200); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6202 = 8'h3a == _T_15 ? $signed(32'sh0) : $signed(_GEN_6201); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6203 = 8'h3b == _T_15 ? $signed(32'sh0) : $signed(_GEN_6202); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6204 = 8'h3c == _T_15 ? $signed(regsB_3_im) : $signed(_GEN_6203); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6205 = 8'h3d == _T_15 ? $signed(regsB_13_im) : $signed(_GEN_6204); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6206 = 8'h3e == _T_15 ? $signed(regsB_23_im) : $signed(_GEN_6205); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6207 = 8'h3f == _T_15 ? $signed(regsB_33_im) : $signed(_GEN_6206); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6208 = 8'h40 == _T_15 ? $signed(regsB_43_im) : $signed(_GEN_6207); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6209 = 8'h41 == _T_15 ? $signed(regsB_53_im) : $signed(_GEN_6208); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6210 = 8'h42 == _T_15 ? $signed(regsB_63_im) : $signed(_GEN_6209); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6211 = 8'h43 == _T_15 ? $signed(regsB_73_im) : $signed(_GEN_6210); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6212 = 8'h44 == _T_15 ? $signed(regsB_83_im) : $signed(_GEN_6211); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6213 = 8'h45 == _T_15 ? $signed(regsB_93_im) : $signed(_GEN_6212); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6214 = 8'h46 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6213); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6215 = 8'h47 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6214); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6216 = 8'h48 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6215); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6217 = 8'h49 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6216); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6218 = 8'h4a == _T_15 ? $signed(32'sh0) : $signed(_GEN_6217); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6219 = 8'h4b == _T_15 ? $signed(32'sh0) : $signed(_GEN_6218); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6220 = 8'h4c == _T_15 ? $signed(32'sh0) : $signed(_GEN_6219); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6221 = 8'h4d == _T_15 ? $signed(32'sh0) : $signed(_GEN_6220); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6222 = 8'h4e == _T_15 ? $signed(32'sh0) : $signed(_GEN_6221); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6223 = 8'h4f == _T_15 ? $signed(32'sh0) : $signed(_GEN_6222); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6224 = 8'h50 == _T_15 ? $signed(regsB_4_im) : $signed(_GEN_6223); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6225 = 8'h51 == _T_15 ? $signed(regsB_14_im) : $signed(_GEN_6224); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6226 = 8'h52 == _T_15 ? $signed(regsB_24_im) : $signed(_GEN_6225); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6227 = 8'h53 == _T_15 ? $signed(regsB_34_im) : $signed(_GEN_6226); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6228 = 8'h54 == _T_15 ? $signed(regsB_44_im) : $signed(_GEN_6227); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6229 = 8'h55 == _T_15 ? $signed(regsB_54_im) : $signed(_GEN_6228); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6230 = 8'h56 == _T_15 ? $signed(regsB_64_im) : $signed(_GEN_6229); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6231 = 8'h57 == _T_15 ? $signed(regsB_74_im) : $signed(_GEN_6230); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6232 = 8'h58 == _T_15 ? $signed(regsB_84_im) : $signed(_GEN_6231); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6233 = 8'h59 == _T_15 ? $signed(regsB_94_im) : $signed(_GEN_6232); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6234 = 8'h5a == _T_15 ? $signed(32'sh0) : $signed(_GEN_6233); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6235 = 8'h5b == _T_15 ? $signed(32'sh0) : $signed(_GEN_6234); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6236 = 8'h5c == _T_15 ? $signed(32'sh0) : $signed(_GEN_6235); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6237 = 8'h5d == _T_15 ? $signed(32'sh0) : $signed(_GEN_6236); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6238 = 8'h5e == _T_15 ? $signed(32'sh0) : $signed(_GEN_6237); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6239 = 8'h5f == _T_15 ? $signed(32'sh0) : $signed(_GEN_6238); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6240 = 8'h60 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6239); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6241 = 8'h61 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6240); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6242 = 8'h62 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6241); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6243 = 8'h63 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6242); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6244 = 8'h64 == _T_15 ? $signed(regsB_5_im) : $signed(_GEN_6243); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6245 = 8'h65 == _T_15 ? $signed(regsB_15_im) : $signed(_GEN_6244); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6246 = 8'h66 == _T_15 ? $signed(regsB_25_im) : $signed(_GEN_6245); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6247 = 8'h67 == _T_15 ? $signed(regsB_35_im) : $signed(_GEN_6246); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6248 = 8'h68 == _T_15 ? $signed(regsB_45_im) : $signed(_GEN_6247); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6249 = 8'h69 == _T_15 ? $signed(regsB_55_im) : $signed(_GEN_6248); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6250 = 8'h6a == _T_15 ? $signed(regsB_65_im) : $signed(_GEN_6249); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6251 = 8'h6b == _T_15 ? $signed(regsB_75_im) : $signed(_GEN_6250); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6252 = 8'h6c == _T_15 ? $signed(regsB_85_im) : $signed(_GEN_6251); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6253 = 8'h6d == _T_15 ? $signed(regsB_95_im) : $signed(_GEN_6252); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6254 = 8'h6e == _T_15 ? $signed(32'sh0) : $signed(_GEN_6253); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6255 = 8'h6f == _T_15 ? $signed(32'sh0) : $signed(_GEN_6254); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6256 = 8'h70 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6255); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6257 = 8'h71 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6256); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6258 = 8'h72 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6257); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6259 = 8'h73 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6258); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6260 = 8'h74 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6259); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6261 = 8'h75 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6260); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6262 = 8'h76 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6261); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6263 = 8'h77 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6262); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6264 = 8'h78 == _T_15 ? $signed(regsB_6_im) : $signed(_GEN_6263); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6265 = 8'h79 == _T_15 ? $signed(regsB_16_im) : $signed(_GEN_6264); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6266 = 8'h7a == _T_15 ? $signed(regsB_26_im) : $signed(_GEN_6265); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6267 = 8'h7b == _T_15 ? $signed(regsB_36_im) : $signed(_GEN_6266); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6268 = 8'h7c == _T_15 ? $signed(regsB_46_im) : $signed(_GEN_6267); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6269 = 8'h7d == _T_15 ? $signed(regsB_56_im) : $signed(_GEN_6268); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6270 = 8'h7e == _T_15 ? $signed(regsB_66_im) : $signed(_GEN_6269); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6271 = 8'h7f == _T_15 ? $signed(regsB_76_im) : $signed(_GEN_6270); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6272 = 8'h80 == _T_15 ? $signed(regsB_86_im) : $signed(_GEN_6271); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6273 = 8'h81 == _T_15 ? $signed(regsB_96_im) : $signed(_GEN_6272); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6274 = 8'h82 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6273); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6275 = 8'h83 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6274); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6276 = 8'h84 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6275); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6277 = 8'h85 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6276); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6278 = 8'h86 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6277); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6279 = 8'h87 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6278); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6280 = 8'h88 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6279); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6281 = 8'h89 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6280); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6282 = 8'h8a == _T_15 ? $signed(32'sh0) : $signed(_GEN_6281); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6283 = 8'h8b == _T_15 ? $signed(32'sh0) : $signed(_GEN_6282); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6284 = 8'h8c == _T_15 ? $signed(regsB_7_im) : $signed(_GEN_6283); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6285 = 8'h8d == _T_15 ? $signed(regsB_17_im) : $signed(_GEN_6284); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6286 = 8'h8e == _T_15 ? $signed(regsB_27_im) : $signed(_GEN_6285); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6287 = 8'h8f == _T_15 ? $signed(regsB_37_im) : $signed(_GEN_6286); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6288 = 8'h90 == _T_15 ? $signed(regsB_47_im) : $signed(_GEN_6287); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6289 = 8'h91 == _T_15 ? $signed(regsB_57_im) : $signed(_GEN_6288); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6290 = 8'h92 == _T_15 ? $signed(regsB_67_im) : $signed(_GEN_6289); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6291 = 8'h93 == _T_15 ? $signed(regsB_77_im) : $signed(_GEN_6290); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6292 = 8'h94 == _T_15 ? $signed(regsB_87_im) : $signed(_GEN_6291); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6293 = 8'h95 == _T_15 ? $signed(regsB_97_im) : $signed(_GEN_6292); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6294 = 8'h96 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6293); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6295 = 8'h97 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6294); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6296 = 8'h98 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6295); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6297 = 8'h99 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6296); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6298 = 8'h9a == _T_15 ? $signed(32'sh0) : $signed(_GEN_6297); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6299 = 8'h9b == _T_15 ? $signed(32'sh0) : $signed(_GEN_6298); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6300 = 8'h9c == _T_15 ? $signed(32'sh0) : $signed(_GEN_6299); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6301 = 8'h9d == _T_15 ? $signed(32'sh0) : $signed(_GEN_6300); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6302 = 8'h9e == _T_15 ? $signed(32'sh0) : $signed(_GEN_6301); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6303 = 8'h9f == _T_15 ? $signed(32'sh0) : $signed(_GEN_6302); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6304 = 8'ha0 == _T_15 ? $signed(regsB_8_im) : $signed(_GEN_6303); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6305 = 8'ha1 == _T_15 ? $signed(regsB_18_im) : $signed(_GEN_6304); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6306 = 8'ha2 == _T_15 ? $signed(regsB_28_im) : $signed(_GEN_6305); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6307 = 8'ha3 == _T_15 ? $signed(regsB_38_im) : $signed(_GEN_6306); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6308 = 8'ha4 == _T_15 ? $signed(regsB_48_im) : $signed(_GEN_6307); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6309 = 8'ha5 == _T_15 ? $signed(regsB_58_im) : $signed(_GEN_6308); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6310 = 8'ha6 == _T_15 ? $signed(regsB_68_im) : $signed(_GEN_6309); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6311 = 8'ha7 == _T_15 ? $signed(regsB_78_im) : $signed(_GEN_6310); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6312 = 8'ha8 == _T_15 ? $signed(regsB_88_im) : $signed(_GEN_6311); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6313 = 8'ha9 == _T_15 ? $signed(regsB_98_im) : $signed(_GEN_6312); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6314 = 8'haa == _T_15 ? $signed(32'sh0) : $signed(_GEN_6313); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6315 = 8'hab == _T_15 ? $signed(32'sh0) : $signed(_GEN_6314); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6316 = 8'hac == _T_15 ? $signed(32'sh0) : $signed(_GEN_6315); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6317 = 8'had == _T_15 ? $signed(32'sh0) : $signed(_GEN_6316); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6318 = 8'hae == _T_15 ? $signed(32'sh0) : $signed(_GEN_6317); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6319 = 8'haf == _T_15 ? $signed(32'sh0) : $signed(_GEN_6318); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6320 = 8'hb0 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6319); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6321 = 8'hb1 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6320); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6322 = 8'hb2 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6321); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6323 = 8'hb3 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6322); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6324 = 8'hb4 == _T_15 ? $signed(regsB_9_im) : $signed(_GEN_6323); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6325 = 8'hb5 == _T_15 ? $signed(regsB_19_im) : $signed(_GEN_6324); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6326 = 8'hb6 == _T_15 ? $signed(regsB_29_im) : $signed(_GEN_6325); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6327 = 8'hb7 == _T_15 ? $signed(regsB_39_im) : $signed(_GEN_6326); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6328 = 8'hb8 == _T_15 ? $signed(regsB_49_im) : $signed(_GEN_6327); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6329 = 8'hb9 == _T_15 ? $signed(regsB_59_im) : $signed(_GEN_6328); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6330 = 8'hba == _T_15 ? $signed(regsB_69_im) : $signed(_GEN_6329); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6331 = 8'hbb == _T_15 ? $signed(regsB_79_im) : $signed(_GEN_6330); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6332 = 8'hbc == _T_15 ? $signed(regsB_89_im) : $signed(_GEN_6331); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6333 = 8'hbd == _T_15 ? $signed(regsB_99_im) : $signed(_GEN_6332); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6335 = 8'h1 == _T_15 ? $signed(regsB_10_re) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6336 = 8'h2 == _T_15 ? $signed(regsB_20_re) : $signed(_GEN_6335); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6337 = 8'h3 == _T_15 ? $signed(regsB_30_re) : $signed(_GEN_6336); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6338 = 8'h4 == _T_15 ? $signed(regsB_40_re) : $signed(_GEN_6337); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6339 = 8'h5 == _T_15 ? $signed(regsB_50_re) : $signed(_GEN_6338); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6340 = 8'h6 == _T_15 ? $signed(regsB_60_re) : $signed(_GEN_6339); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6341 = 8'h7 == _T_15 ? $signed(regsB_70_re) : $signed(_GEN_6340); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6342 = 8'h8 == _T_15 ? $signed(regsB_80_re) : $signed(_GEN_6341); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6343 = 8'h9 == _T_15 ? $signed(regsB_90_re) : $signed(_GEN_6342); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6344 = 8'ha == _T_15 ? $signed(32'sh0) : $signed(_GEN_6343); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6345 = 8'hb == _T_15 ? $signed(32'sh0) : $signed(_GEN_6344); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6346 = 8'hc == _T_15 ? $signed(32'sh0) : $signed(_GEN_6345); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6347 = 8'hd == _T_15 ? $signed(32'sh0) : $signed(_GEN_6346); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6348 = 8'he == _T_15 ? $signed(32'sh0) : $signed(_GEN_6347); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6349 = 8'hf == _T_15 ? $signed(32'sh0) : $signed(_GEN_6348); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6350 = 8'h10 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6349); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6351 = 8'h11 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6350); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6352 = 8'h12 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6351); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6353 = 8'h13 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6352); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6354 = 8'h14 == _T_15 ? $signed(regsB_1_re) : $signed(_GEN_6353); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6355 = 8'h15 == _T_15 ? $signed(regsB_11_re) : $signed(_GEN_6354); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6356 = 8'h16 == _T_15 ? $signed(regsB_21_re) : $signed(_GEN_6355); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6357 = 8'h17 == _T_15 ? $signed(regsB_31_re) : $signed(_GEN_6356); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6358 = 8'h18 == _T_15 ? $signed(regsB_41_re) : $signed(_GEN_6357); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6359 = 8'h19 == _T_15 ? $signed(regsB_51_re) : $signed(_GEN_6358); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6360 = 8'h1a == _T_15 ? $signed(regsB_61_re) : $signed(_GEN_6359); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6361 = 8'h1b == _T_15 ? $signed(regsB_71_re) : $signed(_GEN_6360); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6362 = 8'h1c == _T_15 ? $signed(regsB_81_re) : $signed(_GEN_6361); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6363 = 8'h1d == _T_15 ? $signed(regsB_91_re) : $signed(_GEN_6362); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6364 = 8'h1e == _T_15 ? $signed(32'sh0) : $signed(_GEN_6363); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6365 = 8'h1f == _T_15 ? $signed(32'sh0) : $signed(_GEN_6364); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6366 = 8'h20 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6365); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6367 = 8'h21 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6366); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6368 = 8'h22 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6367); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6369 = 8'h23 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6368); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6370 = 8'h24 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6369); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6371 = 8'h25 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6370); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6372 = 8'h26 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6371); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6373 = 8'h27 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6372); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6374 = 8'h28 == _T_15 ? $signed(regsB_2_re) : $signed(_GEN_6373); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6375 = 8'h29 == _T_15 ? $signed(regsB_12_re) : $signed(_GEN_6374); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6376 = 8'h2a == _T_15 ? $signed(regsB_22_re) : $signed(_GEN_6375); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6377 = 8'h2b == _T_15 ? $signed(regsB_32_re) : $signed(_GEN_6376); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6378 = 8'h2c == _T_15 ? $signed(regsB_42_re) : $signed(_GEN_6377); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6379 = 8'h2d == _T_15 ? $signed(regsB_52_re) : $signed(_GEN_6378); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6380 = 8'h2e == _T_15 ? $signed(regsB_62_re) : $signed(_GEN_6379); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6381 = 8'h2f == _T_15 ? $signed(regsB_72_re) : $signed(_GEN_6380); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6382 = 8'h30 == _T_15 ? $signed(regsB_82_re) : $signed(_GEN_6381); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6383 = 8'h31 == _T_15 ? $signed(regsB_92_re) : $signed(_GEN_6382); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6384 = 8'h32 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6383); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6385 = 8'h33 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6384); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6386 = 8'h34 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6385); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6387 = 8'h35 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6386); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6388 = 8'h36 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6387); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6389 = 8'h37 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6388); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6390 = 8'h38 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6389); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6391 = 8'h39 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6390); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6392 = 8'h3a == _T_15 ? $signed(32'sh0) : $signed(_GEN_6391); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6393 = 8'h3b == _T_15 ? $signed(32'sh0) : $signed(_GEN_6392); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6394 = 8'h3c == _T_15 ? $signed(regsB_3_re) : $signed(_GEN_6393); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6395 = 8'h3d == _T_15 ? $signed(regsB_13_re) : $signed(_GEN_6394); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6396 = 8'h3e == _T_15 ? $signed(regsB_23_re) : $signed(_GEN_6395); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6397 = 8'h3f == _T_15 ? $signed(regsB_33_re) : $signed(_GEN_6396); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6398 = 8'h40 == _T_15 ? $signed(regsB_43_re) : $signed(_GEN_6397); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6399 = 8'h41 == _T_15 ? $signed(regsB_53_re) : $signed(_GEN_6398); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6400 = 8'h42 == _T_15 ? $signed(regsB_63_re) : $signed(_GEN_6399); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6401 = 8'h43 == _T_15 ? $signed(regsB_73_re) : $signed(_GEN_6400); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6402 = 8'h44 == _T_15 ? $signed(regsB_83_re) : $signed(_GEN_6401); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6403 = 8'h45 == _T_15 ? $signed(regsB_93_re) : $signed(_GEN_6402); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6404 = 8'h46 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6403); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6405 = 8'h47 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6404); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6406 = 8'h48 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6405); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6407 = 8'h49 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6406); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6408 = 8'h4a == _T_15 ? $signed(32'sh0) : $signed(_GEN_6407); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6409 = 8'h4b == _T_15 ? $signed(32'sh0) : $signed(_GEN_6408); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6410 = 8'h4c == _T_15 ? $signed(32'sh0) : $signed(_GEN_6409); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6411 = 8'h4d == _T_15 ? $signed(32'sh0) : $signed(_GEN_6410); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6412 = 8'h4e == _T_15 ? $signed(32'sh0) : $signed(_GEN_6411); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6413 = 8'h4f == _T_15 ? $signed(32'sh0) : $signed(_GEN_6412); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6414 = 8'h50 == _T_15 ? $signed(regsB_4_re) : $signed(_GEN_6413); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6415 = 8'h51 == _T_15 ? $signed(regsB_14_re) : $signed(_GEN_6414); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6416 = 8'h52 == _T_15 ? $signed(regsB_24_re) : $signed(_GEN_6415); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6417 = 8'h53 == _T_15 ? $signed(regsB_34_re) : $signed(_GEN_6416); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6418 = 8'h54 == _T_15 ? $signed(regsB_44_re) : $signed(_GEN_6417); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6419 = 8'h55 == _T_15 ? $signed(regsB_54_re) : $signed(_GEN_6418); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6420 = 8'h56 == _T_15 ? $signed(regsB_64_re) : $signed(_GEN_6419); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6421 = 8'h57 == _T_15 ? $signed(regsB_74_re) : $signed(_GEN_6420); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6422 = 8'h58 == _T_15 ? $signed(regsB_84_re) : $signed(_GEN_6421); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6423 = 8'h59 == _T_15 ? $signed(regsB_94_re) : $signed(_GEN_6422); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6424 = 8'h5a == _T_15 ? $signed(32'sh0) : $signed(_GEN_6423); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6425 = 8'h5b == _T_15 ? $signed(32'sh0) : $signed(_GEN_6424); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6426 = 8'h5c == _T_15 ? $signed(32'sh0) : $signed(_GEN_6425); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6427 = 8'h5d == _T_15 ? $signed(32'sh0) : $signed(_GEN_6426); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6428 = 8'h5e == _T_15 ? $signed(32'sh0) : $signed(_GEN_6427); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6429 = 8'h5f == _T_15 ? $signed(32'sh0) : $signed(_GEN_6428); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6430 = 8'h60 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6429); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6431 = 8'h61 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6430); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6432 = 8'h62 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6431); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6433 = 8'h63 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6432); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6434 = 8'h64 == _T_15 ? $signed(regsB_5_re) : $signed(_GEN_6433); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6435 = 8'h65 == _T_15 ? $signed(regsB_15_re) : $signed(_GEN_6434); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6436 = 8'h66 == _T_15 ? $signed(regsB_25_re) : $signed(_GEN_6435); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6437 = 8'h67 == _T_15 ? $signed(regsB_35_re) : $signed(_GEN_6436); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6438 = 8'h68 == _T_15 ? $signed(regsB_45_re) : $signed(_GEN_6437); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6439 = 8'h69 == _T_15 ? $signed(regsB_55_re) : $signed(_GEN_6438); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6440 = 8'h6a == _T_15 ? $signed(regsB_65_re) : $signed(_GEN_6439); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6441 = 8'h6b == _T_15 ? $signed(regsB_75_re) : $signed(_GEN_6440); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6442 = 8'h6c == _T_15 ? $signed(regsB_85_re) : $signed(_GEN_6441); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6443 = 8'h6d == _T_15 ? $signed(regsB_95_re) : $signed(_GEN_6442); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6444 = 8'h6e == _T_15 ? $signed(32'sh0) : $signed(_GEN_6443); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6445 = 8'h6f == _T_15 ? $signed(32'sh0) : $signed(_GEN_6444); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6446 = 8'h70 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6445); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6447 = 8'h71 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6446); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6448 = 8'h72 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6447); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6449 = 8'h73 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6448); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6450 = 8'h74 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6449); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6451 = 8'h75 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6450); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6452 = 8'h76 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6451); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6453 = 8'h77 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6452); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6454 = 8'h78 == _T_15 ? $signed(regsB_6_re) : $signed(_GEN_6453); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6455 = 8'h79 == _T_15 ? $signed(regsB_16_re) : $signed(_GEN_6454); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6456 = 8'h7a == _T_15 ? $signed(regsB_26_re) : $signed(_GEN_6455); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6457 = 8'h7b == _T_15 ? $signed(regsB_36_re) : $signed(_GEN_6456); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6458 = 8'h7c == _T_15 ? $signed(regsB_46_re) : $signed(_GEN_6457); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6459 = 8'h7d == _T_15 ? $signed(regsB_56_re) : $signed(_GEN_6458); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6460 = 8'h7e == _T_15 ? $signed(regsB_66_re) : $signed(_GEN_6459); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6461 = 8'h7f == _T_15 ? $signed(regsB_76_re) : $signed(_GEN_6460); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6462 = 8'h80 == _T_15 ? $signed(regsB_86_re) : $signed(_GEN_6461); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6463 = 8'h81 == _T_15 ? $signed(regsB_96_re) : $signed(_GEN_6462); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6464 = 8'h82 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6463); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6465 = 8'h83 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6464); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6466 = 8'h84 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6465); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6467 = 8'h85 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6466); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6468 = 8'h86 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6467); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6469 = 8'h87 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6468); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6470 = 8'h88 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6469); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6471 = 8'h89 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6470); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6472 = 8'h8a == _T_15 ? $signed(32'sh0) : $signed(_GEN_6471); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6473 = 8'h8b == _T_15 ? $signed(32'sh0) : $signed(_GEN_6472); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6474 = 8'h8c == _T_15 ? $signed(regsB_7_re) : $signed(_GEN_6473); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6475 = 8'h8d == _T_15 ? $signed(regsB_17_re) : $signed(_GEN_6474); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6476 = 8'h8e == _T_15 ? $signed(regsB_27_re) : $signed(_GEN_6475); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6477 = 8'h8f == _T_15 ? $signed(regsB_37_re) : $signed(_GEN_6476); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6478 = 8'h90 == _T_15 ? $signed(regsB_47_re) : $signed(_GEN_6477); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6479 = 8'h91 == _T_15 ? $signed(regsB_57_re) : $signed(_GEN_6478); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6480 = 8'h92 == _T_15 ? $signed(regsB_67_re) : $signed(_GEN_6479); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6481 = 8'h93 == _T_15 ? $signed(regsB_77_re) : $signed(_GEN_6480); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6482 = 8'h94 == _T_15 ? $signed(regsB_87_re) : $signed(_GEN_6481); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6483 = 8'h95 == _T_15 ? $signed(regsB_97_re) : $signed(_GEN_6482); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6484 = 8'h96 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6483); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6485 = 8'h97 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6484); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6486 = 8'h98 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6485); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6487 = 8'h99 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6486); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6488 = 8'h9a == _T_15 ? $signed(32'sh0) : $signed(_GEN_6487); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6489 = 8'h9b == _T_15 ? $signed(32'sh0) : $signed(_GEN_6488); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6490 = 8'h9c == _T_15 ? $signed(32'sh0) : $signed(_GEN_6489); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6491 = 8'h9d == _T_15 ? $signed(32'sh0) : $signed(_GEN_6490); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6492 = 8'h9e == _T_15 ? $signed(32'sh0) : $signed(_GEN_6491); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6493 = 8'h9f == _T_15 ? $signed(32'sh0) : $signed(_GEN_6492); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6494 = 8'ha0 == _T_15 ? $signed(regsB_8_re) : $signed(_GEN_6493); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6495 = 8'ha1 == _T_15 ? $signed(regsB_18_re) : $signed(_GEN_6494); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6496 = 8'ha2 == _T_15 ? $signed(regsB_28_re) : $signed(_GEN_6495); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6497 = 8'ha3 == _T_15 ? $signed(regsB_38_re) : $signed(_GEN_6496); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6498 = 8'ha4 == _T_15 ? $signed(regsB_48_re) : $signed(_GEN_6497); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6499 = 8'ha5 == _T_15 ? $signed(regsB_58_re) : $signed(_GEN_6498); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6500 = 8'ha6 == _T_15 ? $signed(regsB_68_re) : $signed(_GEN_6499); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6501 = 8'ha7 == _T_15 ? $signed(regsB_78_re) : $signed(_GEN_6500); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6502 = 8'ha8 == _T_15 ? $signed(regsB_88_re) : $signed(_GEN_6501); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6503 = 8'ha9 == _T_15 ? $signed(regsB_98_re) : $signed(_GEN_6502); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6504 = 8'haa == _T_15 ? $signed(32'sh0) : $signed(_GEN_6503); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6505 = 8'hab == _T_15 ? $signed(32'sh0) : $signed(_GEN_6504); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6506 = 8'hac == _T_15 ? $signed(32'sh0) : $signed(_GEN_6505); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6507 = 8'had == _T_15 ? $signed(32'sh0) : $signed(_GEN_6506); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6508 = 8'hae == _T_15 ? $signed(32'sh0) : $signed(_GEN_6507); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6509 = 8'haf == _T_15 ? $signed(32'sh0) : $signed(_GEN_6508); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6510 = 8'hb0 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6509); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6511 = 8'hb1 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6510); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6512 = 8'hb2 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6511); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6513 = 8'hb3 == _T_15 ? $signed(32'sh0) : $signed(_GEN_6512); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6514 = 8'hb4 == _T_15 ? $signed(regsB_9_re) : $signed(_GEN_6513); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6515 = 8'hb5 == _T_15 ? $signed(regsB_19_re) : $signed(_GEN_6514); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6516 = 8'hb6 == _T_15 ? $signed(regsB_29_re) : $signed(_GEN_6515); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6517 = 8'hb7 == _T_15 ? $signed(regsB_39_re) : $signed(_GEN_6516); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6518 = 8'hb8 == _T_15 ? $signed(regsB_49_re) : $signed(_GEN_6517); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6519 = 8'hb9 == _T_15 ? $signed(regsB_59_re) : $signed(_GEN_6518); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6520 = 8'hba == _T_15 ? $signed(regsB_69_re) : $signed(_GEN_6519); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6521 = 8'hbb == _T_15 ? $signed(regsB_79_re) : $signed(_GEN_6520); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6522 = 8'hbc == _T_15 ? $signed(regsB_89_re) : $signed(_GEN_6521); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6523 = 8'hbd == _T_15 ? $signed(regsB_99_re) : $signed(_GEN_6522); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6525 = 8'h1 == _T_18 ? $signed(regsB_10_im) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6526 = 8'h2 == _T_18 ? $signed(regsB_20_im) : $signed(_GEN_6525); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6527 = 8'h3 == _T_18 ? $signed(regsB_30_im) : $signed(_GEN_6526); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6528 = 8'h4 == _T_18 ? $signed(regsB_40_im) : $signed(_GEN_6527); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6529 = 8'h5 == _T_18 ? $signed(regsB_50_im) : $signed(_GEN_6528); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6530 = 8'h6 == _T_18 ? $signed(regsB_60_im) : $signed(_GEN_6529); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6531 = 8'h7 == _T_18 ? $signed(regsB_70_im) : $signed(_GEN_6530); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6532 = 8'h8 == _T_18 ? $signed(regsB_80_im) : $signed(_GEN_6531); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6533 = 8'h9 == _T_18 ? $signed(regsB_90_im) : $signed(_GEN_6532); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6534 = 8'ha == _T_18 ? $signed(32'sh0) : $signed(_GEN_6533); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6535 = 8'hb == _T_18 ? $signed(32'sh0) : $signed(_GEN_6534); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6536 = 8'hc == _T_18 ? $signed(32'sh0) : $signed(_GEN_6535); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6537 = 8'hd == _T_18 ? $signed(32'sh0) : $signed(_GEN_6536); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6538 = 8'he == _T_18 ? $signed(32'sh0) : $signed(_GEN_6537); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6539 = 8'hf == _T_18 ? $signed(32'sh0) : $signed(_GEN_6538); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6540 = 8'h10 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6539); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6541 = 8'h11 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6540); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6542 = 8'h12 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6541); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6543 = 8'h13 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6542); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6544 = 8'h14 == _T_18 ? $signed(regsB_1_im) : $signed(_GEN_6543); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6545 = 8'h15 == _T_18 ? $signed(regsB_11_im) : $signed(_GEN_6544); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6546 = 8'h16 == _T_18 ? $signed(regsB_21_im) : $signed(_GEN_6545); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6547 = 8'h17 == _T_18 ? $signed(regsB_31_im) : $signed(_GEN_6546); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6548 = 8'h18 == _T_18 ? $signed(regsB_41_im) : $signed(_GEN_6547); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6549 = 8'h19 == _T_18 ? $signed(regsB_51_im) : $signed(_GEN_6548); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6550 = 8'h1a == _T_18 ? $signed(regsB_61_im) : $signed(_GEN_6549); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6551 = 8'h1b == _T_18 ? $signed(regsB_71_im) : $signed(_GEN_6550); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6552 = 8'h1c == _T_18 ? $signed(regsB_81_im) : $signed(_GEN_6551); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6553 = 8'h1d == _T_18 ? $signed(regsB_91_im) : $signed(_GEN_6552); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6554 = 8'h1e == _T_18 ? $signed(32'sh0) : $signed(_GEN_6553); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6555 = 8'h1f == _T_18 ? $signed(32'sh0) : $signed(_GEN_6554); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6556 = 8'h20 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6555); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6557 = 8'h21 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6556); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6558 = 8'h22 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6557); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6559 = 8'h23 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6558); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6560 = 8'h24 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6559); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6561 = 8'h25 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6560); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6562 = 8'h26 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6561); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6563 = 8'h27 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6562); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6564 = 8'h28 == _T_18 ? $signed(regsB_2_im) : $signed(_GEN_6563); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6565 = 8'h29 == _T_18 ? $signed(regsB_12_im) : $signed(_GEN_6564); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6566 = 8'h2a == _T_18 ? $signed(regsB_22_im) : $signed(_GEN_6565); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6567 = 8'h2b == _T_18 ? $signed(regsB_32_im) : $signed(_GEN_6566); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6568 = 8'h2c == _T_18 ? $signed(regsB_42_im) : $signed(_GEN_6567); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6569 = 8'h2d == _T_18 ? $signed(regsB_52_im) : $signed(_GEN_6568); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6570 = 8'h2e == _T_18 ? $signed(regsB_62_im) : $signed(_GEN_6569); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6571 = 8'h2f == _T_18 ? $signed(regsB_72_im) : $signed(_GEN_6570); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6572 = 8'h30 == _T_18 ? $signed(regsB_82_im) : $signed(_GEN_6571); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6573 = 8'h31 == _T_18 ? $signed(regsB_92_im) : $signed(_GEN_6572); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6574 = 8'h32 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6573); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6575 = 8'h33 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6574); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6576 = 8'h34 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6575); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6577 = 8'h35 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6576); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6578 = 8'h36 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6577); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6579 = 8'h37 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6578); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6580 = 8'h38 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6579); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6581 = 8'h39 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6580); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6582 = 8'h3a == _T_18 ? $signed(32'sh0) : $signed(_GEN_6581); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6583 = 8'h3b == _T_18 ? $signed(32'sh0) : $signed(_GEN_6582); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6584 = 8'h3c == _T_18 ? $signed(regsB_3_im) : $signed(_GEN_6583); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6585 = 8'h3d == _T_18 ? $signed(regsB_13_im) : $signed(_GEN_6584); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6586 = 8'h3e == _T_18 ? $signed(regsB_23_im) : $signed(_GEN_6585); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6587 = 8'h3f == _T_18 ? $signed(regsB_33_im) : $signed(_GEN_6586); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6588 = 8'h40 == _T_18 ? $signed(regsB_43_im) : $signed(_GEN_6587); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6589 = 8'h41 == _T_18 ? $signed(regsB_53_im) : $signed(_GEN_6588); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6590 = 8'h42 == _T_18 ? $signed(regsB_63_im) : $signed(_GEN_6589); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6591 = 8'h43 == _T_18 ? $signed(regsB_73_im) : $signed(_GEN_6590); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6592 = 8'h44 == _T_18 ? $signed(regsB_83_im) : $signed(_GEN_6591); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6593 = 8'h45 == _T_18 ? $signed(regsB_93_im) : $signed(_GEN_6592); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6594 = 8'h46 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6593); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6595 = 8'h47 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6594); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6596 = 8'h48 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6595); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6597 = 8'h49 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6596); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6598 = 8'h4a == _T_18 ? $signed(32'sh0) : $signed(_GEN_6597); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6599 = 8'h4b == _T_18 ? $signed(32'sh0) : $signed(_GEN_6598); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6600 = 8'h4c == _T_18 ? $signed(32'sh0) : $signed(_GEN_6599); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6601 = 8'h4d == _T_18 ? $signed(32'sh0) : $signed(_GEN_6600); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6602 = 8'h4e == _T_18 ? $signed(32'sh0) : $signed(_GEN_6601); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6603 = 8'h4f == _T_18 ? $signed(32'sh0) : $signed(_GEN_6602); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6604 = 8'h50 == _T_18 ? $signed(regsB_4_im) : $signed(_GEN_6603); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6605 = 8'h51 == _T_18 ? $signed(regsB_14_im) : $signed(_GEN_6604); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6606 = 8'h52 == _T_18 ? $signed(regsB_24_im) : $signed(_GEN_6605); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6607 = 8'h53 == _T_18 ? $signed(regsB_34_im) : $signed(_GEN_6606); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6608 = 8'h54 == _T_18 ? $signed(regsB_44_im) : $signed(_GEN_6607); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6609 = 8'h55 == _T_18 ? $signed(regsB_54_im) : $signed(_GEN_6608); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6610 = 8'h56 == _T_18 ? $signed(regsB_64_im) : $signed(_GEN_6609); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6611 = 8'h57 == _T_18 ? $signed(regsB_74_im) : $signed(_GEN_6610); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6612 = 8'h58 == _T_18 ? $signed(regsB_84_im) : $signed(_GEN_6611); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6613 = 8'h59 == _T_18 ? $signed(regsB_94_im) : $signed(_GEN_6612); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6614 = 8'h5a == _T_18 ? $signed(32'sh0) : $signed(_GEN_6613); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6615 = 8'h5b == _T_18 ? $signed(32'sh0) : $signed(_GEN_6614); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6616 = 8'h5c == _T_18 ? $signed(32'sh0) : $signed(_GEN_6615); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6617 = 8'h5d == _T_18 ? $signed(32'sh0) : $signed(_GEN_6616); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6618 = 8'h5e == _T_18 ? $signed(32'sh0) : $signed(_GEN_6617); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6619 = 8'h5f == _T_18 ? $signed(32'sh0) : $signed(_GEN_6618); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6620 = 8'h60 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6619); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6621 = 8'h61 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6620); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6622 = 8'h62 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6621); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6623 = 8'h63 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6622); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6624 = 8'h64 == _T_18 ? $signed(regsB_5_im) : $signed(_GEN_6623); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6625 = 8'h65 == _T_18 ? $signed(regsB_15_im) : $signed(_GEN_6624); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6626 = 8'h66 == _T_18 ? $signed(regsB_25_im) : $signed(_GEN_6625); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6627 = 8'h67 == _T_18 ? $signed(regsB_35_im) : $signed(_GEN_6626); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6628 = 8'h68 == _T_18 ? $signed(regsB_45_im) : $signed(_GEN_6627); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6629 = 8'h69 == _T_18 ? $signed(regsB_55_im) : $signed(_GEN_6628); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6630 = 8'h6a == _T_18 ? $signed(regsB_65_im) : $signed(_GEN_6629); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6631 = 8'h6b == _T_18 ? $signed(regsB_75_im) : $signed(_GEN_6630); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6632 = 8'h6c == _T_18 ? $signed(regsB_85_im) : $signed(_GEN_6631); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6633 = 8'h6d == _T_18 ? $signed(regsB_95_im) : $signed(_GEN_6632); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6634 = 8'h6e == _T_18 ? $signed(32'sh0) : $signed(_GEN_6633); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6635 = 8'h6f == _T_18 ? $signed(32'sh0) : $signed(_GEN_6634); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6636 = 8'h70 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6635); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6637 = 8'h71 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6636); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6638 = 8'h72 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6637); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6639 = 8'h73 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6638); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6640 = 8'h74 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6639); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6641 = 8'h75 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6640); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6642 = 8'h76 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6641); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6643 = 8'h77 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6642); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6644 = 8'h78 == _T_18 ? $signed(regsB_6_im) : $signed(_GEN_6643); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6645 = 8'h79 == _T_18 ? $signed(regsB_16_im) : $signed(_GEN_6644); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6646 = 8'h7a == _T_18 ? $signed(regsB_26_im) : $signed(_GEN_6645); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6647 = 8'h7b == _T_18 ? $signed(regsB_36_im) : $signed(_GEN_6646); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6648 = 8'h7c == _T_18 ? $signed(regsB_46_im) : $signed(_GEN_6647); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6649 = 8'h7d == _T_18 ? $signed(regsB_56_im) : $signed(_GEN_6648); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6650 = 8'h7e == _T_18 ? $signed(regsB_66_im) : $signed(_GEN_6649); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6651 = 8'h7f == _T_18 ? $signed(regsB_76_im) : $signed(_GEN_6650); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6652 = 8'h80 == _T_18 ? $signed(regsB_86_im) : $signed(_GEN_6651); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6653 = 8'h81 == _T_18 ? $signed(regsB_96_im) : $signed(_GEN_6652); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6654 = 8'h82 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6653); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6655 = 8'h83 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6654); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6656 = 8'h84 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6655); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6657 = 8'h85 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6656); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6658 = 8'h86 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6657); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6659 = 8'h87 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6658); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6660 = 8'h88 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6659); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6661 = 8'h89 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6660); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6662 = 8'h8a == _T_18 ? $signed(32'sh0) : $signed(_GEN_6661); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6663 = 8'h8b == _T_18 ? $signed(32'sh0) : $signed(_GEN_6662); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6664 = 8'h8c == _T_18 ? $signed(regsB_7_im) : $signed(_GEN_6663); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6665 = 8'h8d == _T_18 ? $signed(regsB_17_im) : $signed(_GEN_6664); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6666 = 8'h8e == _T_18 ? $signed(regsB_27_im) : $signed(_GEN_6665); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6667 = 8'h8f == _T_18 ? $signed(regsB_37_im) : $signed(_GEN_6666); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6668 = 8'h90 == _T_18 ? $signed(regsB_47_im) : $signed(_GEN_6667); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6669 = 8'h91 == _T_18 ? $signed(regsB_57_im) : $signed(_GEN_6668); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6670 = 8'h92 == _T_18 ? $signed(regsB_67_im) : $signed(_GEN_6669); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6671 = 8'h93 == _T_18 ? $signed(regsB_77_im) : $signed(_GEN_6670); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6672 = 8'h94 == _T_18 ? $signed(regsB_87_im) : $signed(_GEN_6671); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6673 = 8'h95 == _T_18 ? $signed(regsB_97_im) : $signed(_GEN_6672); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6674 = 8'h96 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6673); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6675 = 8'h97 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6674); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6676 = 8'h98 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6675); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6677 = 8'h99 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6676); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6678 = 8'h9a == _T_18 ? $signed(32'sh0) : $signed(_GEN_6677); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6679 = 8'h9b == _T_18 ? $signed(32'sh0) : $signed(_GEN_6678); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6680 = 8'h9c == _T_18 ? $signed(32'sh0) : $signed(_GEN_6679); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6681 = 8'h9d == _T_18 ? $signed(32'sh0) : $signed(_GEN_6680); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6682 = 8'h9e == _T_18 ? $signed(32'sh0) : $signed(_GEN_6681); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6683 = 8'h9f == _T_18 ? $signed(32'sh0) : $signed(_GEN_6682); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6684 = 8'ha0 == _T_18 ? $signed(regsB_8_im) : $signed(_GEN_6683); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6685 = 8'ha1 == _T_18 ? $signed(regsB_18_im) : $signed(_GEN_6684); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6686 = 8'ha2 == _T_18 ? $signed(regsB_28_im) : $signed(_GEN_6685); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6687 = 8'ha3 == _T_18 ? $signed(regsB_38_im) : $signed(_GEN_6686); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6688 = 8'ha4 == _T_18 ? $signed(regsB_48_im) : $signed(_GEN_6687); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6689 = 8'ha5 == _T_18 ? $signed(regsB_58_im) : $signed(_GEN_6688); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6690 = 8'ha6 == _T_18 ? $signed(regsB_68_im) : $signed(_GEN_6689); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6691 = 8'ha7 == _T_18 ? $signed(regsB_78_im) : $signed(_GEN_6690); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6692 = 8'ha8 == _T_18 ? $signed(regsB_88_im) : $signed(_GEN_6691); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6693 = 8'ha9 == _T_18 ? $signed(regsB_98_im) : $signed(_GEN_6692); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6694 = 8'haa == _T_18 ? $signed(32'sh0) : $signed(_GEN_6693); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6695 = 8'hab == _T_18 ? $signed(32'sh0) : $signed(_GEN_6694); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6696 = 8'hac == _T_18 ? $signed(32'sh0) : $signed(_GEN_6695); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6697 = 8'had == _T_18 ? $signed(32'sh0) : $signed(_GEN_6696); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6698 = 8'hae == _T_18 ? $signed(32'sh0) : $signed(_GEN_6697); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6699 = 8'haf == _T_18 ? $signed(32'sh0) : $signed(_GEN_6698); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6700 = 8'hb0 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6699); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6701 = 8'hb1 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6700); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6702 = 8'hb2 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6701); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6703 = 8'hb3 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6702); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6704 = 8'hb4 == _T_18 ? $signed(regsB_9_im) : $signed(_GEN_6703); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6705 = 8'hb5 == _T_18 ? $signed(regsB_19_im) : $signed(_GEN_6704); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6706 = 8'hb6 == _T_18 ? $signed(regsB_29_im) : $signed(_GEN_6705); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6707 = 8'hb7 == _T_18 ? $signed(regsB_39_im) : $signed(_GEN_6706); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6708 = 8'hb8 == _T_18 ? $signed(regsB_49_im) : $signed(_GEN_6707); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6709 = 8'hb9 == _T_18 ? $signed(regsB_59_im) : $signed(_GEN_6708); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6710 = 8'hba == _T_18 ? $signed(regsB_69_im) : $signed(_GEN_6709); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6711 = 8'hbb == _T_18 ? $signed(regsB_79_im) : $signed(_GEN_6710); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6712 = 8'hbc == _T_18 ? $signed(regsB_89_im) : $signed(_GEN_6711); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6713 = 8'hbd == _T_18 ? $signed(regsB_99_im) : $signed(_GEN_6712); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6715 = 8'h1 == _T_18 ? $signed(regsB_10_re) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6716 = 8'h2 == _T_18 ? $signed(regsB_20_re) : $signed(_GEN_6715); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6717 = 8'h3 == _T_18 ? $signed(regsB_30_re) : $signed(_GEN_6716); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6718 = 8'h4 == _T_18 ? $signed(regsB_40_re) : $signed(_GEN_6717); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6719 = 8'h5 == _T_18 ? $signed(regsB_50_re) : $signed(_GEN_6718); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6720 = 8'h6 == _T_18 ? $signed(regsB_60_re) : $signed(_GEN_6719); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6721 = 8'h7 == _T_18 ? $signed(regsB_70_re) : $signed(_GEN_6720); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6722 = 8'h8 == _T_18 ? $signed(regsB_80_re) : $signed(_GEN_6721); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6723 = 8'h9 == _T_18 ? $signed(regsB_90_re) : $signed(_GEN_6722); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6724 = 8'ha == _T_18 ? $signed(32'sh0) : $signed(_GEN_6723); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6725 = 8'hb == _T_18 ? $signed(32'sh0) : $signed(_GEN_6724); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6726 = 8'hc == _T_18 ? $signed(32'sh0) : $signed(_GEN_6725); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6727 = 8'hd == _T_18 ? $signed(32'sh0) : $signed(_GEN_6726); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6728 = 8'he == _T_18 ? $signed(32'sh0) : $signed(_GEN_6727); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6729 = 8'hf == _T_18 ? $signed(32'sh0) : $signed(_GEN_6728); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6730 = 8'h10 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6729); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6731 = 8'h11 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6730); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6732 = 8'h12 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6731); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6733 = 8'h13 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6732); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6734 = 8'h14 == _T_18 ? $signed(regsB_1_re) : $signed(_GEN_6733); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6735 = 8'h15 == _T_18 ? $signed(regsB_11_re) : $signed(_GEN_6734); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6736 = 8'h16 == _T_18 ? $signed(regsB_21_re) : $signed(_GEN_6735); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6737 = 8'h17 == _T_18 ? $signed(regsB_31_re) : $signed(_GEN_6736); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6738 = 8'h18 == _T_18 ? $signed(regsB_41_re) : $signed(_GEN_6737); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6739 = 8'h19 == _T_18 ? $signed(regsB_51_re) : $signed(_GEN_6738); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6740 = 8'h1a == _T_18 ? $signed(regsB_61_re) : $signed(_GEN_6739); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6741 = 8'h1b == _T_18 ? $signed(regsB_71_re) : $signed(_GEN_6740); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6742 = 8'h1c == _T_18 ? $signed(regsB_81_re) : $signed(_GEN_6741); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6743 = 8'h1d == _T_18 ? $signed(regsB_91_re) : $signed(_GEN_6742); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6744 = 8'h1e == _T_18 ? $signed(32'sh0) : $signed(_GEN_6743); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6745 = 8'h1f == _T_18 ? $signed(32'sh0) : $signed(_GEN_6744); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6746 = 8'h20 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6745); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6747 = 8'h21 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6746); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6748 = 8'h22 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6747); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6749 = 8'h23 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6748); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6750 = 8'h24 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6749); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6751 = 8'h25 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6750); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6752 = 8'h26 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6751); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6753 = 8'h27 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6752); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6754 = 8'h28 == _T_18 ? $signed(regsB_2_re) : $signed(_GEN_6753); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6755 = 8'h29 == _T_18 ? $signed(regsB_12_re) : $signed(_GEN_6754); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6756 = 8'h2a == _T_18 ? $signed(regsB_22_re) : $signed(_GEN_6755); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6757 = 8'h2b == _T_18 ? $signed(regsB_32_re) : $signed(_GEN_6756); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6758 = 8'h2c == _T_18 ? $signed(regsB_42_re) : $signed(_GEN_6757); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6759 = 8'h2d == _T_18 ? $signed(regsB_52_re) : $signed(_GEN_6758); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6760 = 8'h2e == _T_18 ? $signed(regsB_62_re) : $signed(_GEN_6759); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6761 = 8'h2f == _T_18 ? $signed(regsB_72_re) : $signed(_GEN_6760); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6762 = 8'h30 == _T_18 ? $signed(regsB_82_re) : $signed(_GEN_6761); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6763 = 8'h31 == _T_18 ? $signed(regsB_92_re) : $signed(_GEN_6762); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6764 = 8'h32 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6763); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6765 = 8'h33 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6764); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6766 = 8'h34 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6765); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6767 = 8'h35 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6766); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6768 = 8'h36 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6767); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6769 = 8'h37 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6768); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6770 = 8'h38 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6769); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6771 = 8'h39 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6770); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6772 = 8'h3a == _T_18 ? $signed(32'sh0) : $signed(_GEN_6771); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6773 = 8'h3b == _T_18 ? $signed(32'sh0) : $signed(_GEN_6772); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6774 = 8'h3c == _T_18 ? $signed(regsB_3_re) : $signed(_GEN_6773); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6775 = 8'h3d == _T_18 ? $signed(regsB_13_re) : $signed(_GEN_6774); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6776 = 8'h3e == _T_18 ? $signed(regsB_23_re) : $signed(_GEN_6775); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6777 = 8'h3f == _T_18 ? $signed(regsB_33_re) : $signed(_GEN_6776); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6778 = 8'h40 == _T_18 ? $signed(regsB_43_re) : $signed(_GEN_6777); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6779 = 8'h41 == _T_18 ? $signed(regsB_53_re) : $signed(_GEN_6778); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6780 = 8'h42 == _T_18 ? $signed(regsB_63_re) : $signed(_GEN_6779); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6781 = 8'h43 == _T_18 ? $signed(regsB_73_re) : $signed(_GEN_6780); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6782 = 8'h44 == _T_18 ? $signed(regsB_83_re) : $signed(_GEN_6781); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6783 = 8'h45 == _T_18 ? $signed(regsB_93_re) : $signed(_GEN_6782); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6784 = 8'h46 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6783); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6785 = 8'h47 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6784); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6786 = 8'h48 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6785); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6787 = 8'h49 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6786); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6788 = 8'h4a == _T_18 ? $signed(32'sh0) : $signed(_GEN_6787); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6789 = 8'h4b == _T_18 ? $signed(32'sh0) : $signed(_GEN_6788); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6790 = 8'h4c == _T_18 ? $signed(32'sh0) : $signed(_GEN_6789); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6791 = 8'h4d == _T_18 ? $signed(32'sh0) : $signed(_GEN_6790); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6792 = 8'h4e == _T_18 ? $signed(32'sh0) : $signed(_GEN_6791); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6793 = 8'h4f == _T_18 ? $signed(32'sh0) : $signed(_GEN_6792); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6794 = 8'h50 == _T_18 ? $signed(regsB_4_re) : $signed(_GEN_6793); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6795 = 8'h51 == _T_18 ? $signed(regsB_14_re) : $signed(_GEN_6794); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6796 = 8'h52 == _T_18 ? $signed(regsB_24_re) : $signed(_GEN_6795); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6797 = 8'h53 == _T_18 ? $signed(regsB_34_re) : $signed(_GEN_6796); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6798 = 8'h54 == _T_18 ? $signed(regsB_44_re) : $signed(_GEN_6797); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6799 = 8'h55 == _T_18 ? $signed(regsB_54_re) : $signed(_GEN_6798); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6800 = 8'h56 == _T_18 ? $signed(regsB_64_re) : $signed(_GEN_6799); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6801 = 8'h57 == _T_18 ? $signed(regsB_74_re) : $signed(_GEN_6800); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6802 = 8'h58 == _T_18 ? $signed(regsB_84_re) : $signed(_GEN_6801); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6803 = 8'h59 == _T_18 ? $signed(regsB_94_re) : $signed(_GEN_6802); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6804 = 8'h5a == _T_18 ? $signed(32'sh0) : $signed(_GEN_6803); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6805 = 8'h5b == _T_18 ? $signed(32'sh0) : $signed(_GEN_6804); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6806 = 8'h5c == _T_18 ? $signed(32'sh0) : $signed(_GEN_6805); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6807 = 8'h5d == _T_18 ? $signed(32'sh0) : $signed(_GEN_6806); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6808 = 8'h5e == _T_18 ? $signed(32'sh0) : $signed(_GEN_6807); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6809 = 8'h5f == _T_18 ? $signed(32'sh0) : $signed(_GEN_6808); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6810 = 8'h60 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6809); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6811 = 8'h61 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6810); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6812 = 8'h62 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6811); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6813 = 8'h63 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6812); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6814 = 8'h64 == _T_18 ? $signed(regsB_5_re) : $signed(_GEN_6813); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6815 = 8'h65 == _T_18 ? $signed(regsB_15_re) : $signed(_GEN_6814); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6816 = 8'h66 == _T_18 ? $signed(regsB_25_re) : $signed(_GEN_6815); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6817 = 8'h67 == _T_18 ? $signed(regsB_35_re) : $signed(_GEN_6816); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6818 = 8'h68 == _T_18 ? $signed(regsB_45_re) : $signed(_GEN_6817); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6819 = 8'h69 == _T_18 ? $signed(regsB_55_re) : $signed(_GEN_6818); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6820 = 8'h6a == _T_18 ? $signed(regsB_65_re) : $signed(_GEN_6819); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6821 = 8'h6b == _T_18 ? $signed(regsB_75_re) : $signed(_GEN_6820); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6822 = 8'h6c == _T_18 ? $signed(regsB_85_re) : $signed(_GEN_6821); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6823 = 8'h6d == _T_18 ? $signed(regsB_95_re) : $signed(_GEN_6822); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6824 = 8'h6e == _T_18 ? $signed(32'sh0) : $signed(_GEN_6823); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6825 = 8'h6f == _T_18 ? $signed(32'sh0) : $signed(_GEN_6824); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6826 = 8'h70 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6825); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6827 = 8'h71 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6826); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6828 = 8'h72 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6827); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6829 = 8'h73 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6828); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6830 = 8'h74 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6829); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6831 = 8'h75 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6830); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6832 = 8'h76 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6831); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6833 = 8'h77 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6832); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6834 = 8'h78 == _T_18 ? $signed(regsB_6_re) : $signed(_GEN_6833); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6835 = 8'h79 == _T_18 ? $signed(regsB_16_re) : $signed(_GEN_6834); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6836 = 8'h7a == _T_18 ? $signed(regsB_26_re) : $signed(_GEN_6835); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6837 = 8'h7b == _T_18 ? $signed(regsB_36_re) : $signed(_GEN_6836); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6838 = 8'h7c == _T_18 ? $signed(regsB_46_re) : $signed(_GEN_6837); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6839 = 8'h7d == _T_18 ? $signed(regsB_56_re) : $signed(_GEN_6838); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6840 = 8'h7e == _T_18 ? $signed(regsB_66_re) : $signed(_GEN_6839); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6841 = 8'h7f == _T_18 ? $signed(regsB_76_re) : $signed(_GEN_6840); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6842 = 8'h80 == _T_18 ? $signed(regsB_86_re) : $signed(_GEN_6841); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6843 = 8'h81 == _T_18 ? $signed(regsB_96_re) : $signed(_GEN_6842); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6844 = 8'h82 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6843); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6845 = 8'h83 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6844); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6846 = 8'h84 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6845); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6847 = 8'h85 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6846); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6848 = 8'h86 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6847); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6849 = 8'h87 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6848); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6850 = 8'h88 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6849); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6851 = 8'h89 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6850); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6852 = 8'h8a == _T_18 ? $signed(32'sh0) : $signed(_GEN_6851); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6853 = 8'h8b == _T_18 ? $signed(32'sh0) : $signed(_GEN_6852); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6854 = 8'h8c == _T_18 ? $signed(regsB_7_re) : $signed(_GEN_6853); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6855 = 8'h8d == _T_18 ? $signed(regsB_17_re) : $signed(_GEN_6854); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6856 = 8'h8e == _T_18 ? $signed(regsB_27_re) : $signed(_GEN_6855); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6857 = 8'h8f == _T_18 ? $signed(regsB_37_re) : $signed(_GEN_6856); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6858 = 8'h90 == _T_18 ? $signed(regsB_47_re) : $signed(_GEN_6857); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6859 = 8'h91 == _T_18 ? $signed(regsB_57_re) : $signed(_GEN_6858); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6860 = 8'h92 == _T_18 ? $signed(regsB_67_re) : $signed(_GEN_6859); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6861 = 8'h93 == _T_18 ? $signed(regsB_77_re) : $signed(_GEN_6860); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6862 = 8'h94 == _T_18 ? $signed(regsB_87_re) : $signed(_GEN_6861); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6863 = 8'h95 == _T_18 ? $signed(regsB_97_re) : $signed(_GEN_6862); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6864 = 8'h96 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6863); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6865 = 8'h97 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6864); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6866 = 8'h98 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6865); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6867 = 8'h99 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6866); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6868 = 8'h9a == _T_18 ? $signed(32'sh0) : $signed(_GEN_6867); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6869 = 8'h9b == _T_18 ? $signed(32'sh0) : $signed(_GEN_6868); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6870 = 8'h9c == _T_18 ? $signed(32'sh0) : $signed(_GEN_6869); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6871 = 8'h9d == _T_18 ? $signed(32'sh0) : $signed(_GEN_6870); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6872 = 8'h9e == _T_18 ? $signed(32'sh0) : $signed(_GEN_6871); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6873 = 8'h9f == _T_18 ? $signed(32'sh0) : $signed(_GEN_6872); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6874 = 8'ha0 == _T_18 ? $signed(regsB_8_re) : $signed(_GEN_6873); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6875 = 8'ha1 == _T_18 ? $signed(regsB_18_re) : $signed(_GEN_6874); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6876 = 8'ha2 == _T_18 ? $signed(regsB_28_re) : $signed(_GEN_6875); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6877 = 8'ha3 == _T_18 ? $signed(regsB_38_re) : $signed(_GEN_6876); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6878 = 8'ha4 == _T_18 ? $signed(regsB_48_re) : $signed(_GEN_6877); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6879 = 8'ha5 == _T_18 ? $signed(regsB_58_re) : $signed(_GEN_6878); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6880 = 8'ha6 == _T_18 ? $signed(regsB_68_re) : $signed(_GEN_6879); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6881 = 8'ha7 == _T_18 ? $signed(regsB_78_re) : $signed(_GEN_6880); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6882 = 8'ha8 == _T_18 ? $signed(regsB_88_re) : $signed(_GEN_6881); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6883 = 8'ha9 == _T_18 ? $signed(regsB_98_re) : $signed(_GEN_6882); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6884 = 8'haa == _T_18 ? $signed(32'sh0) : $signed(_GEN_6883); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6885 = 8'hab == _T_18 ? $signed(32'sh0) : $signed(_GEN_6884); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6886 = 8'hac == _T_18 ? $signed(32'sh0) : $signed(_GEN_6885); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6887 = 8'had == _T_18 ? $signed(32'sh0) : $signed(_GEN_6886); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6888 = 8'hae == _T_18 ? $signed(32'sh0) : $signed(_GEN_6887); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6889 = 8'haf == _T_18 ? $signed(32'sh0) : $signed(_GEN_6888); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6890 = 8'hb0 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6889); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6891 = 8'hb1 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6890); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6892 = 8'hb2 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6891); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6893 = 8'hb3 == _T_18 ? $signed(32'sh0) : $signed(_GEN_6892); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6894 = 8'hb4 == _T_18 ? $signed(regsB_9_re) : $signed(_GEN_6893); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6895 = 8'hb5 == _T_18 ? $signed(regsB_19_re) : $signed(_GEN_6894); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6896 = 8'hb6 == _T_18 ? $signed(regsB_29_re) : $signed(_GEN_6895); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6897 = 8'hb7 == _T_18 ? $signed(regsB_39_re) : $signed(_GEN_6896); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6898 = 8'hb8 == _T_18 ? $signed(regsB_49_re) : $signed(_GEN_6897); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6899 = 8'hb9 == _T_18 ? $signed(regsB_59_re) : $signed(_GEN_6898); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6900 = 8'hba == _T_18 ? $signed(regsB_69_re) : $signed(_GEN_6899); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6901 = 8'hbb == _T_18 ? $signed(regsB_79_re) : $signed(_GEN_6900); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6902 = 8'hbc == _T_18 ? $signed(regsB_89_re) : $signed(_GEN_6901); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6903 = 8'hbd == _T_18 ? $signed(regsB_99_re) : $signed(_GEN_6902); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6905 = 8'h1 == _T_21 ? $signed(regsB_10_im) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6906 = 8'h2 == _T_21 ? $signed(regsB_20_im) : $signed(_GEN_6905); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6907 = 8'h3 == _T_21 ? $signed(regsB_30_im) : $signed(_GEN_6906); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6908 = 8'h4 == _T_21 ? $signed(regsB_40_im) : $signed(_GEN_6907); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6909 = 8'h5 == _T_21 ? $signed(regsB_50_im) : $signed(_GEN_6908); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6910 = 8'h6 == _T_21 ? $signed(regsB_60_im) : $signed(_GEN_6909); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6911 = 8'h7 == _T_21 ? $signed(regsB_70_im) : $signed(_GEN_6910); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6912 = 8'h8 == _T_21 ? $signed(regsB_80_im) : $signed(_GEN_6911); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6913 = 8'h9 == _T_21 ? $signed(regsB_90_im) : $signed(_GEN_6912); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6914 = 8'ha == _T_21 ? $signed(32'sh0) : $signed(_GEN_6913); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6915 = 8'hb == _T_21 ? $signed(32'sh0) : $signed(_GEN_6914); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6916 = 8'hc == _T_21 ? $signed(32'sh0) : $signed(_GEN_6915); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6917 = 8'hd == _T_21 ? $signed(32'sh0) : $signed(_GEN_6916); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6918 = 8'he == _T_21 ? $signed(32'sh0) : $signed(_GEN_6917); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6919 = 8'hf == _T_21 ? $signed(32'sh0) : $signed(_GEN_6918); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6920 = 8'h10 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6919); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6921 = 8'h11 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6920); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6922 = 8'h12 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6921); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6923 = 8'h13 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6922); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6924 = 8'h14 == _T_21 ? $signed(regsB_1_im) : $signed(_GEN_6923); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6925 = 8'h15 == _T_21 ? $signed(regsB_11_im) : $signed(_GEN_6924); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6926 = 8'h16 == _T_21 ? $signed(regsB_21_im) : $signed(_GEN_6925); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6927 = 8'h17 == _T_21 ? $signed(regsB_31_im) : $signed(_GEN_6926); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6928 = 8'h18 == _T_21 ? $signed(regsB_41_im) : $signed(_GEN_6927); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6929 = 8'h19 == _T_21 ? $signed(regsB_51_im) : $signed(_GEN_6928); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6930 = 8'h1a == _T_21 ? $signed(regsB_61_im) : $signed(_GEN_6929); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6931 = 8'h1b == _T_21 ? $signed(regsB_71_im) : $signed(_GEN_6930); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6932 = 8'h1c == _T_21 ? $signed(regsB_81_im) : $signed(_GEN_6931); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6933 = 8'h1d == _T_21 ? $signed(regsB_91_im) : $signed(_GEN_6932); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6934 = 8'h1e == _T_21 ? $signed(32'sh0) : $signed(_GEN_6933); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6935 = 8'h1f == _T_21 ? $signed(32'sh0) : $signed(_GEN_6934); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6936 = 8'h20 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6935); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6937 = 8'h21 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6936); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6938 = 8'h22 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6937); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6939 = 8'h23 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6938); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6940 = 8'h24 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6939); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6941 = 8'h25 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6940); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6942 = 8'h26 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6941); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6943 = 8'h27 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6942); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6944 = 8'h28 == _T_21 ? $signed(regsB_2_im) : $signed(_GEN_6943); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6945 = 8'h29 == _T_21 ? $signed(regsB_12_im) : $signed(_GEN_6944); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6946 = 8'h2a == _T_21 ? $signed(regsB_22_im) : $signed(_GEN_6945); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6947 = 8'h2b == _T_21 ? $signed(regsB_32_im) : $signed(_GEN_6946); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6948 = 8'h2c == _T_21 ? $signed(regsB_42_im) : $signed(_GEN_6947); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6949 = 8'h2d == _T_21 ? $signed(regsB_52_im) : $signed(_GEN_6948); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6950 = 8'h2e == _T_21 ? $signed(regsB_62_im) : $signed(_GEN_6949); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6951 = 8'h2f == _T_21 ? $signed(regsB_72_im) : $signed(_GEN_6950); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6952 = 8'h30 == _T_21 ? $signed(regsB_82_im) : $signed(_GEN_6951); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6953 = 8'h31 == _T_21 ? $signed(regsB_92_im) : $signed(_GEN_6952); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6954 = 8'h32 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6953); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6955 = 8'h33 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6954); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6956 = 8'h34 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6955); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6957 = 8'h35 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6956); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6958 = 8'h36 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6957); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6959 = 8'h37 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6958); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6960 = 8'h38 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6959); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6961 = 8'h39 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6960); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6962 = 8'h3a == _T_21 ? $signed(32'sh0) : $signed(_GEN_6961); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6963 = 8'h3b == _T_21 ? $signed(32'sh0) : $signed(_GEN_6962); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6964 = 8'h3c == _T_21 ? $signed(regsB_3_im) : $signed(_GEN_6963); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6965 = 8'h3d == _T_21 ? $signed(regsB_13_im) : $signed(_GEN_6964); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6966 = 8'h3e == _T_21 ? $signed(regsB_23_im) : $signed(_GEN_6965); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6967 = 8'h3f == _T_21 ? $signed(regsB_33_im) : $signed(_GEN_6966); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6968 = 8'h40 == _T_21 ? $signed(regsB_43_im) : $signed(_GEN_6967); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6969 = 8'h41 == _T_21 ? $signed(regsB_53_im) : $signed(_GEN_6968); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6970 = 8'h42 == _T_21 ? $signed(regsB_63_im) : $signed(_GEN_6969); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6971 = 8'h43 == _T_21 ? $signed(regsB_73_im) : $signed(_GEN_6970); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6972 = 8'h44 == _T_21 ? $signed(regsB_83_im) : $signed(_GEN_6971); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6973 = 8'h45 == _T_21 ? $signed(regsB_93_im) : $signed(_GEN_6972); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6974 = 8'h46 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6973); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6975 = 8'h47 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6974); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6976 = 8'h48 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6975); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6977 = 8'h49 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6976); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6978 = 8'h4a == _T_21 ? $signed(32'sh0) : $signed(_GEN_6977); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6979 = 8'h4b == _T_21 ? $signed(32'sh0) : $signed(_GEN_6978); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6980 = 8'h4c == _T_21 ? $signed(32'sh0) : $signed(_GEN_6979); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6981 = 8'h4d == _T_21 ? $signed(32'sh0) : $signed(_GEN_6980); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6982 = 8'h4e == _T_21 ? $signed(32'sh0) : $signed(_GEN_6981); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6983 = 8'h4f == _T_21 ? $signed(32'sh0) : $signed(_GEN_6982); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6984 = 8'h50 == _T_21 ? $signed(regsB_4_im) : $signed(_GEN_6983); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6985 = 8'h51 == _T_21 ? $signed(regsB_14_im) : $signed(_GEN_6984); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6986 = 8'h52 == _T_21 ? $signed(regsB_24_im) : $signed(_GEN_6985); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6987 = 8'h53 == _T_21 ? $signed(regsB_34_im) : $signed(_GEN_6986); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6988 = 8'h54 == _T_21 ? $signed(regsB_44_im) : $signed(_GEN_6987); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6989 = 8'h55 == _T_21 ? $signed(regsB_54_im) : $signed(_GEN_6988); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6990 = 8'h56 == _T_21 ? $signed(regsB_64_im) : $signed(_GEN_6989); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6991 = 8'h57 == _T_21 ? $signed(regsB_74_im) : $signed(_GEN_6990); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6992 = 8'h58 == _T_21 ? $signed(regsB_84_im) : $signed(_GEN_6991); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6993 = 8'h59 == _T_21 ? $signed(regsB_94_im) : $signed(_GEN_6992); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6994 = 8'h5a == _T_21 ? $signed(32'sh0) : $signed(_GEN_6993); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6995 = 8'h5b == _T_21 ? $signed(32'sh0) : $signed(_GEN_6994); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6996 = 8'h5c == _T_21 ? $signed(32'sh0) : $signed(_GEN_6995); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6997 = 8'h5d == _T_21 ? $signed(32'sh0) : $signed(_GEN_6996); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6998 = 8'h5e == _T_21 ? $signed(32'sh0) : $signed(_GEN_6997); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_6999 = 8'h5f == _T_21 ? $signed(32'sh0) : $signed(_GEN_6998); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7000 = 8'h60 == _T_21 ? $signed(32'sh0) : $signed(_GEN_6999); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7001 = 8'h61 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7000); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7002 = 8'h62 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7001); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7003 = 8'h63 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7002); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7004 = 8'h64 == _T_21 ? $signed(regsB_5_im) : $signed(_GEN_7003); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7005 = 8'h65 == _T_21 ? $signed(regsB_15_im) : $signed(_GEN_7004); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7006 = 8'h66 == _T_21 ? $signed(regsB_25_im) : $signed(_GEN_7005); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7007 = 8'h67 == _T_21 ? $signed(regsB_35_im) : $signed(_GEN_7006); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7008 = 8'h68 == _T_21 ? $signed(regsB_45_im) : $signed(_GEN_7007); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7009 = 8'h69 == _T_21 ? $signed(regsB_55_im) : $signed(_GEN_7008); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7010 = 8'h6a == _T_21 ? $signed(regsB_65_im) : $signed(_GEN_7009); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7011 = 8'h6b == _T_21 ? $signed(regsB_75_im) : $signed(_GEN_7010); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7012 = 8'h6c == _T_21 ? $signed(regsB_85_im) : $signed(_GEN_7011); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7013 = 8'h6d == _T_21 ? $signed(regsB_95_im) : $signed(_GEN_7012); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7014 = 8'h6e == _T_21 ? $signed(32'sh0) : $signed(_GEN_7013); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7015 = 8'h6f == _T_21 ? $signed(32'sh0) : $signed(_GEN_7014); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7016 = 8'h70 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7015); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7017 = 8'h71 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7016); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7018 = 8'h72 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7017); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7019 = 8'h73 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7018); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7020 = 8'h74 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7019); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7021 = 8'h75 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7020); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7022 = 8'h76 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7021); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7023 = 8'h77 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7022); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7024 = 8'h78 == _T_21 ? $signed(regsB_6_im) : $signed(_GEN_7023); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7025 = 8'h79 == _T_21 ? $signed(regsB_16_im) : $signed(_GEN_7024); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7026 = 8'h7a == _T_21 ? $signed(regsB_26_im) : $signed(_GEN_7025); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7027 = 8'h7b == _T_21 ? $signed(regsB_36_im) : $signed(_GEN_7026); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7028 = 8'h7c == _T_21 ? $signed(regsB_46_im) : $signed(_GEN_7027); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7029 = 8'h7d == _T_21 ? $signed(regsB_56_im) : $signed(_GEN_7028); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7030 = 8'h7e == _T_21 ? $signed(regsB_66_im) : $signed(_GEN_7029); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7031 = 8'h7f == _T_21 ? $signed(regsB_76_im) : $signed(_GEN_7030); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7032 = 8'h80 == _T_21 ? $signed(regsB_86_im) : $signed(_GEN_7031); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7033 = 8'h81 == _T_21 ? $signed(regsB_96_im) : $signed(_GEN_7032); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7034 = 8'h82 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7033); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7035 = 8'h83 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7034); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7036 = 8'h84 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7035); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7037 = 8'h85 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7036); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7038 = 8'h86 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7037); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7039 = 8'h87 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7038); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7040 = 8'h88 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7039); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7041 = 8'h89 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7040); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7042 = 8'h8a == _T_21 ? $signed(32'sh0) : $signed(_GEN_7041); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7043 = 8'h8b == _T_21 ? $signed(32'sh0) : $signed(_GEN_7042); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7044 = 8'h8c == _T_21 ? $signed(regsB_7_im) : $signed(_GEN_7043); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7045 = 8'h8d == _T_21 ? $signed(regsB_17_im) : $signed(_GEN_7044); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7046 = 8'h8e == _T_21 ? $signed(regsB_27_im) : $signed(_GEN_7045); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7047 = 8'h8f == _T_21 ? $signed(regsB_37_im) : $signed(_GEN_7046); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7048 = 8'h90 == _T_21 ? $signed(regsB_47_im) : $signed(_GEN_7047); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7049 = 8'h91 == _T_21 ? $signed(regsB_57_im) : $signed(_GEN_7048); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7050 = 8'h92 == _T_21 ? $signed(regsB_67_im) : $signed(_GEN_7049); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7051 = 8'h93 == _T_21 ? $signed(regsB_77_im) : $signed(_GEN_7050); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7052 = 8'h94 == _T_21 ? $signed(regsB_87_im) : $signed(_GEN_7051); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7053 = 8'h95 == _T_21 ? $signed(regsB_97_im) : $signed(_GEN_7052); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7054 = 8'h96 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7053); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7055 = 8'h97 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7054); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7056 = 8'h98 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7055); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7057 = 8'h99 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7056); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7058 = 8'h9a == _T_21 ? $signed(32'sh0) : $signed(_GEN_7057); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7059 = 8'h9b == _T_21 ? $signed(32'sh0) : $signed(_GEN_7058); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7060 = 8'h9c == _T_21 ? $signed(32'sh0) : $signed(_GEN_7059); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7061 = 8'h9d == _T_21 ? $signed(32'sh0) : $signed(_GEN_7060); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7062 = 8'h9e == _T_21 ? $signed(32'sh0) : $signed(_GEN_7061); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7063 = 8'h9f == _T_21 ? $signed(32'sh0) : $signed(_GEN_7062); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7064 = 8'ha0 == _T_21 ? $signed(regsB_8_im) : $signed(_GEN_7063); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7065 = 8'ha1 == _T_21 ? $signed(regsB_18_im) : $signed(_GEN_7064); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7066 = 8'ha2 == _T_21 ? $signed(regsB_28_im) : $signed(_GEN_7065); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7067 = 8'ha3 == _T_21 ? $signed(regsB_38_im) : $signed(_GEN_7066); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7068 = 8'ha4 == _T_21 ? $signed(regsB_48_im) : $signed(_GEN_7067); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7069 = 8'ha5 == _T_21 ? $signed(regsB_58_im) : $signed(_GEN_7068); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7070 = 8'ha6 == _T_21 ? $signed(regsB_68_im) : $signed(_GEN_7069); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7071 = 8'ha7 == _T_21 ? $signed(regsB_78_im) : $signed(_GEN_7070); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7072 = 8'ha8 == _T_21 ? $signed(regsB_88_im) : $signed(_GEN_7071); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7073 = 8'ha9 == _T_21 ? $signed(regsB_98_im) : $signed(_GEN_7072); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7074 = 8'haa == _T_21 ? $signed(32'sh0) : $signed(_GEN_7073); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7075 = 8'hab == _T_21 ? $signed(32'sh0) : $signed(_GEN_7074); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7076 = 8'hac == _T_21 ? $signed(32'sh0) : $signed(_GEN_7075); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7077 = 8'had == _T_21 ? $signed(32'sh0) : $signed(_GEN_7076); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7078 = 8'hae == _T_21 ? $signed(32'sh0) : $signed(_GEN_7077); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7079 = 8'haf == _T_21 ? $signed(32'sh0) : $signed(_GEN_7078); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7080 = 8'hb0 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7079); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7081 = 8'hb1 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7080); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7082 = 8'hb2 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7081); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7083 = 8'hb3 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7082); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7084 = 8'hb4 == _T_21 ? $signed(regsB_9_im) : $signed(_GEN_7083); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7085 = 8'hb5 == _T_21 ? $signed(regsB_19_im) : $signed(_GEN_7084); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7086 = 8'hb6 == _T_21 ? $signed(regsB_29_im) : $signed(_GEN_7085); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7087 = 8'hb7 == _T_21 ? $signed(regsB_39_im) : $signed(_GEN_7086); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7088 = 8'hb8 == _T_21 ? $signed(regsB_49_im) : $signed(_GEN_7087); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7089 = 8'hb9 == _T_21 ? $signed(regsB_59_im) : $signed(_GEN_7088); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7090 = 8'hba == _T_21 ? $signed(regsB_69_im) : $signed(_GEN_7089); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7091 = 8'hbb == _T_21 ? $signed(regsB_79_im) : $signed(_GEN_7090); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7092 = 8'hbc == _T_21 ? $signed(regsB_89_im) : $signed(_GEN_7091); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7093 = 8'hbd == _T_21 ? $signed(regsB_99_im) : $signed(_GEN_7092); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7095 = 8'h1 == _T_21 ? $signed(regsB_10_re) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7096 = 8'h2 == _T_21 ? $signed(regsB_20_re) : $signed(_GEN_7095); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7097 = 8'h3 == _T_21 ? $signed(regsB_30_re) : $signed(_GEN_7096); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7098 = 8'h4 == _T_21 ? $signed(regsB_40_re) : $signed(_GEN_7097); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7099 = 8'h5 == _T_21 ? $signed(regsB_50_re) : $signed(_GEN_7098); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7100 = 8'h6 == _T_21 ? $signed(regsB_60_re) : $signed(_GEN_7099); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7101 = 8'h7 == _T_21 ? $signed(regsB_70_re) : $signed(_GEN_7100); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7102 = 8'h8 == _T_21 ? $signed(regsB_80_re) : $signed(_GEN_7101); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7103 = 8'h9 == _T_21 ? $signed(regsB_90_re) : $signed(_GEN_7102); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7104 = 8'ha == _T_21 ? $signed(32'sh0) : $signed(_GEN_7103); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7105 = 8'hb == _T_21 ? $signed(32'sh0) : $signed(_GEN_7104); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7106 = 8'hc == _T_21 ? $signed(32'sh0) : $signed(_GEN_7105); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7107 = 8'hd == _T_21 ? $signed(32'sh0) : $signed(_GEN_7106); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7108 = 8'he == _T_21 ? $signed(32'sh0) : $signed(_GEN_7107); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7109 = 8'hf == _T_21 ? $signed(32'sh0) : $signed(_GEN_7108); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7110 = 8'h10 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7109); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7111 = 8'h11 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7110); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7112 = 8'h12 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7111); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7113 = 8'h13 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7112); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7114 = 8'h14 == _T_21 ? $signed(regsB_1_re) : $signed(_GEN_7113); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7115 = 8'h15 == _T_21 ? $signed(regsB_11_re) : $signed(_GEN_7114); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7116 = 8'h16 == _T_21 ? $signed(regsB_21_re) : $signed(_GEN_7115); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7117 = 8'h17 == _T_21 ? $signed(regsB_31_re) : $signed(_GEN_7116); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7118 = 8'h18 == _T_21 ? $signed(regsB_41_re) : $signed(_GEN_7117); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7119 = 8'h19 == _T_21 ? $signed(regsB_51_re) : $signed(_GEN_7118); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7120 = 8'h1a == _T_21 ? $signed(regsB_61_re) : $signed(_GEN_7119); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7121 = 8'h1b == _T_21 ? $signed(regsB_71_re) : $signed(_GEN_7120); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7122 = 8'h1c == _T_21 ? $signed(regsB_81_re) : $signed(_GEN_7121); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7123 = 8'h1d == _T_21 ? $signed(regsB_91_re) : $signed(_GEN_7122); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7124 = 8'h1e == _T_21 ? $signed(32'sh0) : $signed(_GEN_7123); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7125 = 8'h1f == _T_21 ? $signed(32'sh0) : $signed(_GEN_7124); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7126 = 8'h20 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7125); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7127 = 8'h21 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7126); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7128 = 8'h22 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7127); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7129 = 8'h23 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7128); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7130 = 8'h24 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7129); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7131 = 8'h25 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7130); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7132 = 8'h26 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7131); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7133 = 8'h27 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7132); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7134 = 8'h28 == _T_21 ? $signed(regsB_2_re) : $signed(_GEN_7133); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7135 = 8'h29 == _T_21 ? $signed(regsB_12_re) : $signed(_GEN_7134); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7136 = 8'h2a == _T_21 ? $signed(regsB_22_re) : $signed(_GEN_7135); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7137 = 8'h2b == _T_21 ? $signed(regsB_32_re) : $signed(_GEN_7136); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7138 = 8'h2c == _T_21 ? $signed(regsB_42_re) : $signed(_GEN_7137); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7139 = 8'h2d == _T_21 ? $signed(regsB_52_re) : $signed(_GEN_7138); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7140 = 8'h2e == _T_21 ? $signed(regsB_62_re) : $signed(_GEN_7139); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7141 = 8'h2f == _T_21 ? $signed(regsB_72_re) : $signed(_GEN_7140); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7142 = 8'h30 == _T_21 ? $signed(regsB_82_re) : $signed(_GEN_7141); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7143 = 8'h31 == _T_21 ? $signed(regsB_92_re) : $signed(_GEN_7142); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7144 = 8'h32 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7143); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7145 = 8'h33 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7144); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7146 = 8'h34 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7145); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7147 = 8'h35 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7146); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7148 = 8'h36 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7147); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7149 = 8'h37 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7148); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7150 = 8'h38 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7149); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7151 = 8'h39 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7150); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7152 = 8'h3a == _T_21 ? $signed(32'sh0) : $signed(_GEN_7151); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7153 = 8'h3b == _T_21 ? $signed(32'sh0) : $signed(_GEN_7152); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7154 = 8'h3c == _T_21 ? $signed(regsB_3_re) : $signed(_GEN_7153); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7155 = 8'h3d == _T_21 ? $signed(regsB_13_re) : $signed(_GEN_7154); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7156 = 8'h3e == _T_21 ? $signed(regsB_23_re) : $signed(_GEN_7155); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7157 = 8'h3f == _T_21 ? $signed(regsB_33_re) : $signed(_GEN_7156); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7158 = 8'h40 == _T_21 ? $signed(regsB_43_re) : $signed(_GEN_7157); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7159 = 8'h41 == _T_21 ? $signed(regsB_53_re) : $signed(_GEN_7158); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7160 = 8'h42 == _T_21 ? $signed(regsB_63_re) : $signed(_GEN_7159); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7161 = 8'h43 == _T_21 ? $signed(regsB_73_re) : $signed(_GEN_7160); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7162 = 8'h44 == _T_21 ? $signed(regsB_83_re) : $signed(_GEN_7161); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7163 = 8'h45 == _T_21 ? $signed(regsB_93_re) : $signed(_GEN_7162); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7164 = 8'h46 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7163); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7165 = 8'h47 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7164); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7166 = 8'h48 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7165); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7167 = 8'h49 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7166); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7168 = 8'h4a == _T_21 ? $signed(32'sh0) : $signed(_GEN_7167); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7169 = 8'h4b == _T_21 ? $signed(32'sh0) : $signed(_GEN_7168); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7170 = 8'h4c == _T_21 ? $signed(32'sh0) : $signed(_GEN_7169); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7171 = 8'h4d == _T_21 ? $signed(32'sh0) : $signed(_GEN_7170); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7172 = 8'h4e == _T_21 ? $signed(32'sh0) : $signed(_GEN_7171); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7173 = 8'h4f == _T_21 ? $signed(32'sh0) : $signed(_GEN_7172); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7174 = 8'h50 == _T_21 ? $signed(regsB_4_re) : $signed(_GEN_7173); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7175 = 8'h51 == _T_21 ? $signed(regsB_14_re) : $signed(_GEN_7174); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7176 = 8'h52 == _T_21 ? $signed(regsB_24_re) : $signed(_GEN_7175); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7177 = 8'h53 == _T_21 ? $signed(regsB_34_re) : $signed(_GEN_7176); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7178 = 8'h54 == _T_21 ? $signed(regsB_44_re) : $signed(_GEN_7177); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7179 = 8'h55 == _T_21 ? $signed(regsB_54_re) : $signed(_GEN_7178); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7180 = 8'h56 == _T_21 ? $signed(regsB_64_re) : $signed(_GEN_7179); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7181 = 8'h57 == _T_21 ? $signed(regsB_74_re) : $signed(_GEN_7180); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7182 = 8'h58 == _T_21 ? $signed(regsB_84_re) : $signed(_GEN_7181); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7183 = 8'h59 == _T_21 ? $signed(regsB_94_re) : $signed(_GEN_7182); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7184 = 8'h5a == _T_21 ? $signed(32'sh0) : $signed(_GEN_7183); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7185 = 8'h5b == _T_21 ? $signed(32'sh0) : $signed(_GEN_7184); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7186 = 8'h5c == _T_21 ? $signed(32'sh0) : $signed(_GEN_7185); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7187 = 8'h5d == _T_21 ? $signed(32'sh0) : $signed(_GEN_7186); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7188 = 8'h5e == _T_21 ? $signed(32'sh0) : $signed(_GEN_7187); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7189 = 8'h5f == _T_21 ? $signed(32'sh0) : $signed(_GEN_7188); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7190 = 8'h60 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7189); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7191 = 8'h61 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7190); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7192 = 8'h62 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7191); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7193 = 8'h63 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7192); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7194 = 8'h64 == _T_21 ? $signed(regsB_5_re) : $signed(_GEN_7193); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7195 = 8'h65 == _T_21 ? $signed(regsB_15_re) : $signed(_GEN_7194); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7196 = 8'h66 == _T_21 ? $signed(regsB_25_re) : $signed(_GEN_7195); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7197 = 8'h67 == _T_21 ? $signed(regsB_35_re) : $signed(_GEN_7196); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7198 = 8'h68 == _T_21 ? $signed(regsB_45_re) : $signed(_GEN_7197); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7199 = 8'h69 == _T_21 ? $signed(regsB_55_re) : $signed(_GEN_7198); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7200 = 8'h6a == _T_21 ? $signed(regsB_65_re) : $signed(_GEN_7199); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7201 = 8'h6b == _T_21 ? $signed(regsB_75_re) : $signed(_GEN_7200); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7202 = 8'h6c == _T_21 ? $signed(regsB_85_re) : $signed(_GEN_7201); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7203 = 8'h6d == _T_21 ? $signed(regsB_95_re) : $signed(_GEN_7202); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7204 = 8'h6e == _T_21 ? $signed(32'sh0) : $signed(_GEN_7203); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7205 = 8'h6f == _T_21 ? $signed(32'sh0) : $signed(_GEN_7204); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7206 = 8'h70 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7205); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7207 = 8'h71 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7206); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7208 = 8'h72 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7207); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7209 = 8'h73 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7208); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7210 = 8'h74 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7209); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7211 = 8'h75 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7210); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7212 = 8'h76 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7211); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7213 = 8'h77 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7212); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7214 = 8'h78 == _T_21 ? $signed(regsB_6_re) : $signed(_GEN_7213); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7215 = 8'h79 == _T_21 ? $signed(regsB_16_re) : $signed(_GEN_7214); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7216 = 8'h7a == _T_21 ? $signed(regsB_26_re) : $signed(_GEN_7215); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7217 = 8'h7b == _T_21 ? $signed(regsB_36_re) : $signed(_GEN_7216); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7218 = 8'h7c == _T_21 ? $signed(regsB_46_re) : $signed(_GEN_7217); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7219 = 8'h7d == _T_21 ? $signed(regsB_56_re) : $signed(_GEN_7218); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7220 = 8'h7e == _T_21 ? $signed(regsB_66_re) : $signed(_GEN_7219); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7221 = 8'h7f == _T_21 ? $signed(regsB_76_re) : $signed(_GEN_7220); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7222 = 8'h80 == _T_21 ? $signed(regsB_86_re) : $signed(_GEN_7221); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7223 = 8'h81 == _T_21 ? $signed(regsB_96_re) : $signed(_GEN_7222); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7224 = 8'h82 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7223); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7225 = 8'h83 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7224); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7226 = 8'h84 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7225); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7227 = 8'h85 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7226); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7228 = 8'h86 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7227); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7229 = 8'h87 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7228); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7230 = 8'h88 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7229); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7231 = 8'h89 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7230); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7232 = 8'h8a == _T_21 ? $signed(32'sh0) : $signed(_GEN_7231); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7233 = 8'h8b == _T_21 ? $signed(32'sh0) : $signed(_GEN_7232); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7234 = 8'h8c == _T_21 ? $signed(regsB_7_re) : $signed(_GEN_7233); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7235 = 8'h8d == _T_21 ? $signed(regsB_17_re) : $signed(_GEN_7234); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7236 = 8'h8e == _T_21 ? $signed(regsB_27_re) : $signed(_GEN_7235); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7237 = 8'h8f == _T_21 ? $signed(regsB_37_re) : $signed(_GEN_7236); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7238 = 8'h90 == _T_21 ? $signed(regsB_47_re) : $signed(_GEN_7237); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7239 = 8'h91 == _T_21 ? $signed(regsB_57_re) : $signed(_GEN_7238); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7240 = 8'h92 == _T_21 ? $signed(regsB_67_re) : $signed(_GEN_7239); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7241 = 8'h93 == _T_21 ? $signed(regsB_77_re) : $signed(_GEN_7240); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7242 = 8'h94 == _T_21 ? $signed(regsB_87_re) : $signed(_GEN_7241); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7243 = 8'h95 == _T_21 ? $signed(regsB_97_re) : $signed(_GEN_7242); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7244 = 8'h96 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7243); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7245 = 8'h97 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7244); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7246 = 8'h98 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7245); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7247 = 8'h99 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7246); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7248 = 8'h9a == _T_21 ? $signed(32'sh0) : $signed(_GEN_7247); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7249 = 8'h9b == _T_21 ? $signed(32'sh0) : $signed(_GEN_7248); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7250 = 8'h9c == _T_21 ? $signed(32'sh0) : $signed(_GEN_7249); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7251 = 8'h9d == _T_21 ? $signed(32'sh0) : $signed(_GEN_7250); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7252 = 8'h9e == _T_21 ? $signed(32'sh0) : $signed(_GEN_7251); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7253 = 8'h9f == _T_21 ? $signed(32'sh0) : $signed(_GEN_7252); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7254 = 8'ha0 == _T_21 ? $signed(regsB_8_re) : $signed(_GEN_7253); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7255 = 8'ha1 == _T_21 ? $signed(regsB_18_re) : $signed(_GEN_7254); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7256 = 8'ha2 == _T_21 ? $signed(regsB_28_re) : $signed(_GEN_7255); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7257 = 8'ha3 == _T_21 ? $signed(regsB_38_re) : $signed(_GEN_7256); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7258 = 8'ha4 == _T_21 ? $signed(regsB_48_re) : $signed(_GEN_7257); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7259 = 8'ha5 == _T_21 ? $signed(regsB_58_re) : $signed(_GEN_7258); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7260 = 8'ha6 == _T_21 ? $signed(regsB_68_re) : $signed(_GEN_7259); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7261 = 8'ha7 == _T_21 ? $signed(regsB_78_re) : $signed(_GEN_7260); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7262 = 8'ha8 == _T_21 ? $signed(regsB_88_re) : $signed(_GEN_7261); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7263 = 8'ha9 == _T_21 ? $signed(regsB_98_re) : $signed(_GEN_7262); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7264 = 8'haa == _T_21 ? $signed(32'sh0) : $signed(_GEN_7263); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7265 = 8'hab == _T_21 ? $signed(32'sh0) : $signed(_GEN_7264); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7266 = 8'hac == _T_21 ? $signed(32'sh0) : $signed(_GEN_7265); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7267 = 8'had == _T_21 ? $signed(32'sh0) : $signed(_GEN_7266); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7268 = 8'hae == _T_21 ? $signed(32'sh0) : $signed(_GEN_7267); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7269 = 8'haf == _T_21 ? $signed(32'sh0) : $signed(_GEN_7268); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7270 = 8'hb0 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7269); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7271 = 8'hb1 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7270); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7272 = 8'hb2 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7271); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7273 = 8'hb3 == _T_21 ? $signed(32'sh0) : $signed(_GEN_7272); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7274 = 8'hb4 == _T_21 ? $signed(regsB_9_re) : $signed(_GEN_7273); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7275 = 8'hb5 == _T_21 ? $signed(regsB_19_re) : $signed(_GEN_7274); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7276 = 8'hb6 == _T_21 ? $signed(regsB_29_re) : $signed(_GEN_7275); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7277 = 8'hb7 == _T_21 ? $signed(regsB_39_re) : $signed(_GEN_7276); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7278 = 8'hb8 == _T_21 ? $signed(regsB_49_re) : $signed(_GEN_7277); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7279 = 8'hb9 == _T_21 ? $signed(regsB_59_re) : $signed(_GEN_7278); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7280 = 8'hba == _T_21 ? $signed(regsB_69_re) : $signed(_GEN_7279); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7281 = 8'hbb == _T_21 ? $signed(regsB_79_re) : $signed(_GEN_7280); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7282 = 8'hbc == _T_21 ? $signed(regsB_89_re) : $signed(_GEN_7281); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7283 = 8'hbd == _T_21 ? $signed(regsB_99_re) : $signed(_GEN_7282); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7285 = 8'h1 == _T_24 ? $signed(regsB_10_im) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7286 = 8'h2 == _T_24 ? $signed(regsB_20_im) : $signed(_GEN_7285); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7287 = 8'h3 == _T_24 ? $signed(regsB_30_im) : $signed(_GEN_7286); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7288 = 8'h4 == _T_24 ? $signed(regsB_40_im) : $signed(_GEN_7287); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7289 = 8'h5 == _T_24 ? $signed(regsB_50_im) : $signed(_GEN_7288); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7290 = 8'h6 == _T_24 ? $signed(regsB_60_im) : $signed(_GEN_7289); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7291 = 8'h7 == _T_24 ? $signed(regsB_70_im) : $signed(_GEN_7290); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7292 = 8'h8 == _T_24 ? $signed(regsB_80_im) : $signed(_GEN_7291); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7293 = 8'h9 == _T_24 ? $signed(regsB_90_im) : $signed(_GEN_7292); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7294 = 8'ha == _T_24 ? $signed(32'sh0) : $signed(_GEN_7293); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7295 = 8'hb == _T_24 ? $signed(32'sh0) : $signed(_GEN_7294); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7296 = 8'hc == _T_24 ? $signed(32'sh0) : $signed(_GEN_7295); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7297 = 8'hd == _T_24 ? $signed(32'sh0) : $signed(_GEN_7296); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7298 = 8'he == _T_24 ? $signed(32'sh0) : $signed(_GEN_7297); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7299 = 8'hf == _T_24 ? $signed(32'sh0) : $signed(_GEN_7298); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7300 = 8'h10 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7299); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7301 = 8'h11 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7300); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7302 = 8'h12 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7301); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7303 = 8'h13 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7302); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7304 = 8'h14 == _T_24 ? $signed(regsB_1_im) : $signed(_GEN_7303); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7305 = 8'h15 == _T_24 ? $signed(regsB_11_im) : $signed(_GEN_7304); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7306 = 8'h16 == _T_24 ? $signed(regsB_21_im) : $signed(_GEN_7305); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7307 = 8'h17 == _T_24 ? $signed(regsB_31_im) : $signed(_GEN_7306); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7308 = 8'h18 == _T_24 ? $signed(regsB_41_im) : $signed(_GEN_7307); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7309 = 8'h19 == _T_24 ? $signed(regsB_51_im) : $signed(_GEN_7308); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7310 = 8'h1a == _T_24 ? $signed(regsB_61_im) : $signed(_GEN_7309); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7311 = 8'h1b == _T_24 ? $signed(regsB_71_im) : $signed(_GEN_7310); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7312 = 8'h1c == _T_24 ? $signed(regsB_81_im) : $signed(_GEN_7311); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7313 = 8'h1d == _T_24 ? $signed(regsB_91_im) : $signed(_GEN_7312); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7314 = 8'h1e == _T_24 ? $signed(32'sh0) : $signed(_GEN_7313); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7315 = 8'h1f == _T_24 ? $signed(32'sh0) : $signed(_GEN_7314); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7316 = 8'h20 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7315); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7317 = 8'h21 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7316); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7318 = 8'h22 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7317); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7319 = 8'h23 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7318); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7320 = 8'h24 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7319); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7321 = 8'h25 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7320); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7322 = 8'h26 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7321); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7323 = 8'h27 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7322); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7324 = 8'h28 == _T_24 ? $signed(regsB_2_im) : $signed(_GEN_7323); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7325 = 8'h29 == _T_24 ? $signed(regsB_12_im) : $signed(_GEN_7324); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7326 = 8'h2a == _T_24 ? $signed(regsB_22_im) : $signed(_GEN_7325); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7327 = 8'h2b == _T_24 ? $signed(regsB_32_im) : $signed(_GEN_7326); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7328 = 8'h2c == _T_24 ? $signed(regsB_42_im) : $signed(_GEN_7327); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7329 = 8'h2d == _T_24 ? $signed(regsB_52_im) : $signed(_GEN_7328); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7330 = 8'h2e == _T_24 ? $signed(regsB_62_im) : $signed(_GEN_7329); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7331 = 8'h2f == _T_24 ? $signed(regsB_72_im) : $signed(_GEN_7330); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7332 = 8'h30 == _T_24 ? $signed(regsB_82_im) : $signed(_GEN_7331); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7333 = 8'h31 == _T_24 ? $signed(regsB_92_im) : $signed(_GEN_7332); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7334 = 8'h32 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7333); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7335 = 8'h33 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7334); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7336 = 8'h34 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7335); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7337 = 8'h35 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7336); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7338 = 8'h36 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7337); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7339 = 8'h37 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7338); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7340 = 8'h38 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7339); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7341 = 8'h39 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7340); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7342 = 8'h3a == _T_24 ? $signed(32'sh0) : $signed(_GEN_7341); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7343 = 8'h3b == _T_24 ? $signed(32'sh0) : $signed(_GEN_7342); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7344 = 8'h3c == _T_24 ? $signed(regsB_3_im) : $signed(_GEN_7343); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7345 = 8'h3d == _T_24 ? $signed(regsB_13_im) : $signed(_GEN_7344); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7346 = 8'h3e == _T_24 ? $signed(regsB_23_im) : $signed(_GEN_7345); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7347 = 8'h3f == _T_24 ? $signed(regsB_33_im) : $signed(_GEN_7346); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7348 = 8'h40 == _T_24 ? $signed(regsB_43_im) : $signed(_GEN_7347); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7349 = 8'h41 == _T_24 ? $signed(regsB_53_im) : $signed(_GEN_7348); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7350 = 8'h42 == _T_24 ? $signed(regsB_63_im) : $signed(_GEN_7349); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7351 = 8'h43 == _T_24 ? $signed(regsB_73_im) : $signed(_GEN_7350); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7352 = 8'h44 == _T_24 ? $signed(regsB_83_im) : $signed(_GEN_7351); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7353 = 8'h45 == _T_24 ? $signed(regsB_93_im) : $signed(_GEN_7352); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7354 = 8'h46 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7353); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7355 = 8'h47 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7354); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7356 = 8'h48 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7355); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7357 = 8'h49 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7356); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7358 = 8'h4a == _T_24 ? $signed(32'sh0) : $signed(_GEN_7357); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7359 = 8'h4b == _T_24 ? $signed(32'sh0) : $signed(_GEN_7358); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7360 = 8'h4c == _T_24 ? $signed(32'sh0) : $signed(_GEN_7359); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7361 = 8'h4d == _T_24 ? $signed(32'sh0) : $signed(_GEN_7360); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7362 = 8'h4e == _T_24 ? $signed(32'sh0) : $signed(_GEN_7361); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7363 = 8'h4f == _T_24 ? $signed(32'sh0) : $signed(_GEN_7362); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7364 = 8'h50 == _T_24 ? $signed(regsB_4_im) : $signed(_GEN_7363); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7365 = 8'h51 == _T_24 ? $signed(regsB_14_im) : $signed(_GEN_7364); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7366 = 8'h52 == _T_24 ? $signed(regsB_24_im) : $signed(_GEN_7365); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7367 = 8'h53 == _T_24 ? $signed(regsB_34_im) : $signed(_GEN_7366); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7368 = 8'h54 == _T_24 ? $signed(regsB_44_im) : $signed(_GEN_7367); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7369 = 8'h55 == _T_24 ? $signed(regsB_54_im) : $signed(_GEN_7368); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7370 = 8'h56 == _T_24 ? $signed(regsB_64_im) : $signed(_GEN_7369); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7371 = 8'h57 == _T_24 ? $signed(regsB_74_im) : $signed(_GEN_7370); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7372 = 8'h58 == _T_24 ? $signed(regsB_84_im) : $signed(_GEN_7371); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7373 = 8'h59 == _T_24 ? $signed(regsB_94_im) : $signed(_GEN_7372); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7374 = 8'h5a == _T_24 ? $signed(32'sh0) : $signed(_GEN_7373); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7375 = 8'h5b == _T_24 ? $signed(32'sh0) : $signed(_GEN_7374); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7376 = 8'h5c == _T_24 ? $signed(32'sh0) : $signed(_GEN_7375); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7377 = 8'h5d == _T_24 ? $signed(32'sh0) : $signed(_GEN_7376); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7378 = 8'h5e == _T_24 ? $signed(32'sh0) : $signed(_GEN_7377); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7379 = 8'h5f == _T_24 ? $signed(32'sh0) : $signed(_GEN_7378); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7380 = 8'h60 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7379); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7381 = 8'h61 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7380); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7382 = 8'h62 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7381); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7383 = 8'h63 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7382); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7384 = 8'h64 == _T_24 ? $signed(regsB_5_im) : $signed(_GEN_7383); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7385 = 8'h65 == _T_24 ? $signed(regsB_15_im) : $signed(_GEN_7384); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7386 = 8'h66 == _T_24 ? $signed(regsB_25_im) : $signed(_GEN_7385); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7387 = 8'h67 == _T_24 ? $signed(regsB_35_im) : $signed(_GEN_7386); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7388 = 8'h68 == _T_24 ? $signed(regsB_45_im) : $signed(_GEN_7387); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7389 = 8'h69 == _T_24 ? $signed(regsB_55_im) : $signed(_GEN_7388); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7390 = 8'h6a == _T_24 ? $signed(regsB_65_im) : $signed(_GEN_7389); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7391 = 8'h6b == _T_24 ? $signed(regsB_75_im) : $signed(_GEN_7390); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7392 = 8'h6c == _T_24 ? $signed(regsB_85_im) : $signed(_GEN_7391); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7393 = 8'h6d == _T_24 ? $signed(regsB_95_im) : $signed(_GEN_7392); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7394 = 8'h6e == _T_24 ? $signed(32'sh0) : $signed(_GEN_7393); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7395 = 8'h6f == _T_24 ? $signed(32'sh0) : $signed(_GEN_7394); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7396 = 8'h70 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7395); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7397 = 8'h71 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7396); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7398 = 8'h72 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7397); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7399 = 8'h73 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7398); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7400 = 8'h74 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7399); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7401 = 8'h75 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7400); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7402 = 8'h76 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7401); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7403 = 8'h77 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7402); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7404 = 8'h78 == _T_24 ? $signed(regsB_6_im) : $signed(_GEN_7403); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7405 = 8'h79 == _T_24 ? $signed(regsB_16_im) : $signed(_GEN_7404); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7406 = 8'h7a == _T_24 ? $signed(regsB_26_im) : $signed(_GEN_7405); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7407 = 8'h7b == _T_24 ? $signed(regsB_36_im) : $signed(_GEN_7406); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7408 = 8'h7c == _T_24 ? $signed(regsB_46_im) : $signed(_GEN_7407); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7409 = 8'h7d == _T_24 ? $signed(regsB_56_im) : $signed(_GEN_7408); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7410 = 8'h7e == _T_24 ? $signed(regsB_66_im) : $signed(_GEN_7409); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7411 = 8'h7f == _T_24 ? $signed(regsB_76_im) : $signed(_GEN_7410); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7412 = 8'h80 == _T_24 ? $signed(regsB_86_im) : $signed(_GEN_7411); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7413 = 8'h81 == _T_24 ? $signed(regsB_96_im) : $signed(_GEN_7412); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7414 = 8'h82 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7413); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7415 = 8'h83 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7414); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7416 = 8'h84 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7415); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7417 = 8'h85 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7416); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7418 = 8'h86 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7417); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7419 = 8'h87 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7418); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7420 = 8'h88 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7419); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7421 = 8'h89 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7420); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7422 = 8'h8a == _T_24 ? $signed(32'sh0) : $signed(_GEN_7421); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7423 = 8'h8b == _T_24 ? $signed(32'sh0) : $signed(_GEN_7422); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7424 = 8'h8c == _T_24 ? $signed(regsB_7_im) : $signed(_GEN_7423); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7425 = 8'h8d == _T_24 ? $signed(regsB_17_im) : $signed(_GEN_7424); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7426 = 8'h8e == _T_24 ? $signed(regsB_27_im) : $signed(_GEN_7425); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7427 = 8'h8f == _T_24 ? $signed(regsB_37_im) : $signed(_GEN_7426); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7428 = 8'h90 == _T_24 ? $signed(regsB_47_im) : $signed(_GEN_7427); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7429 = 8'h91 == _T_24 ? $signed(regsB_57_im) : $signed(_GEN_7428); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7430 = 8'h92 == _T_24 ? $signed(regsB_67_im) : $signed(_GEN_7429); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7431 = 8'h93 == _T_24 ? $signed(regsB_77_im) : $signed(_GEN_7430); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7432 = 8'h94 == _T_24 ? $signed(regsB_87_im) : $signed(_GEN_7431); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7433 = 8'h95 == _T_24 ? $signed(regsB_97_im) : $signed(_GEN_7432); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7434 = 8'h96 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7433); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7435 = 8'h97 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7434); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7436 = 8'h98 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7435); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7437 = 8'h99 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7436); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7438 = 8'h9a == _T_24 ? $signed(32'sh0) : $signed(_GEN_7437); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7439 = 8'h9b == _T_24 ? $signed(32'sh0) : $signed(_GEN_7438); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7440 = 8'h9c == _T_24 ? $signed(32'sh0) : $signed(_GEN_7439); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7441 = 8'h9d == _T_24 ? $signed(32'sh0) : $signed(_GEN_7440); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7442 = 8'h9e == _T_24 ? $signed(32'sh0) : $signed(_GEN_7441); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7443 = 8'h9f == _T_24 ? $signed(32'sh0) : $signed(_GEN_7442); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7444 = 8'ha0 == _T_24 ? $signed(regsB_8_im) : $signed(_GEN_7443); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7445 = 8'ha1 == _T_24 ? $signed(regsB_18_im) : $signed(_GEN_7444); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7446 = 8'ha2 == _T_24 ? $signed(regsB_28_im) : $signed(_GEN_7445); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7447 = 8'ha3 == _T_24 ? $signed(regsB_38_im) : $signed(_GEN_7446); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7448 = 8'ha4 == _T_24 ? $signed(regsB_48_im) : $signed(_GEN_7447); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7449 = 8'ha5 == _T_24 ? $signed(regsB_58_im) : $signed(_GEN_7448); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7450 = 8'ha6 == _T_24 ? $signed(regsB_68_im) : $signed(_GEN_7449); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7451 = 8'ha7 == _T_24 ? $signed(regsB_78_im) : $signed(_GEN_7450); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7452 = 8'ha8 == _T_24 ? $signed(regsB_88_im) : $signed(_GEN_7451); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7453 = 8'ha9 == _T_24 ? $signed(regsB_98_im) : $signed(_GEN_7452); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7454 = 8'haa == _T_24 ? $signed(32'sh0) : $signed(_GEN_7453); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7455 = 8'hab == _T_24 ? $signed(32'sh0) : $signed(_GEN_7454); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7456 = 8'hac == _T_24 ? $signed(32'sh0) : $signed(_GEN_7455); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7457 = 8'had == _T_24 ? $signed(32'sh0) : $signed(_GEN_7456); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7458 = 8'hae == _T_24 ? $signed(32'sh0) : $signed(_GEN_7457); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7459 = 8'haf == _T_24 ? $signed(32'sh0) : $signed(_GEN_7458); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7460 = 8'hb0 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7459); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7461 = 8'hb1 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7460); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7462 = 8'hb2 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7461); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7463 = 8'hb3 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7462); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7464 = 8'hb4 == _T_24 ? $signed(regsB_9_im) : $signed(_GEN_7463); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7465 = 8'hb5 == _T_24 ? $signed(regsB_19_im) : $signed(_GEN_7464); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7466 = 8'hb6 == _T_24 ? $signed(regsB_29_im) : $signed(_GEN_7465); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7467 = 8'hb7 == _T_24 ? $signed(regsB_39_im) : $signed(_GEN_7466); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7468 = 8'hb8 == _T_24 ? $signed(regsB_49_im) : $signed(_GEN_7467); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7469 = 8'hb9 == _T_24 ? $signed(regsB_59_im) : $signed(_GEN_7468); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7470 = 8'hba == _T_24 ? $signed(regsB_69_im) : $signed(_GEN_7469); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7471 = 8'hbb == _T_24 ? $signed(regsB_79_im) : $signed(_GEN_7470); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7472 = 8'hbc == _T_24 ? $signed(regsB_89_im) : $signed(_GEN_7471); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7473 = 8'hbd == _T_24 ? $signed(regsB_99_im) : $signed(_GEN_7472); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7475 = 8'h1 == _T_24 ? $signed(regsB_10_re) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7476 = 8'h2 == _T_24 ? $signed(regsB_20_re) : $signed(_GEN_7475); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7477 = 8'h3 == _T_24 ? $signed(regsB_30_re) : $signed(_GEN_7476); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7478 = 8'h4 == _T_24 ? $signed(regsB_40_re) : $signed(_GEN_7477); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7479 = 8'h5 == _T_24 ? $signed(regsB_50_re) : $signed(_GEN_7478); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7480 = 8'h6 == _T_24 ? $signed(regsB_60_re) : $signed(_GEN_7479); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7481 = 8'h7 == _T_24 ? $signed(regsB_70_re) : $signed(_GEN_7480); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7482 = 8'h8 == _T_24 ? $signed(regsB_80_re) : $signed(_GEN_7481); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7483 = 8'h9 == _T_24 ? $signed(regsB_90_re) : $signed(_GEN_7482); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7484 = 8'ha == _T_24 ? $signed(32'sh0) : $signed(_GEN_7483); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7485 = 8'hb == _T_24 ? $signed(32'sh0) : $signed(_GEN_7484); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7486 = 8'hc == _T_24 ? $signed(32'sh0) : $signed(_GEN_7485); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7487 = 8'hd == _T_24 ? $signed(32'sh0) : $signed(_GEN_7486); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7488 = 8'he == _T_24 ? $signed(32'sh0) : $signed(_GEN_7487); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7489 = 8'hf == _T_24 ? $signed(32'sh0) : $signed(_GEN_7488); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7490 = 8'h10 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7489); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7491 = 8'h11 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7490); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7492 = 8'h12 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7491); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7493 = 8'h13 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7492); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7494 = 8'h14 == _T_24 ? $signed(regsB_1_re) : $signed(_GEN_7493); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7495 = 8'h15 == _T_24 ? $signed(regsB_11_re) : $signed(_GEN_7494); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7496 = 8'h16 == _T_24 ? $signed(regsB_21_re) : $signed(_GEN_7495); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7497 = 8'h17 == _T_24 ? $signed(regsB_31_re) : $signed(_GEN_7496); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7498 = 8'h18 == _T_24 ? $signed(regsB_41_re) : $signed(_GEN_7497); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7499 = 8'h19 == _T_24 ? $signed(regsB_51_re) : $signed(_GEN_7498); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7500 = 8'h1a == _T_24 ? $signed(regsB_61_re) : $signed(_GEN_7499); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7501 = 8'h1b == _T_24 ? $signed(regsB_71_re) : $signed(_GEN_7500); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7502 = 8'h1c == _T_24 ? $signed(regsB_81_re) : $signed(_GEN_7501); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7503 = 8'h1d == _T_24 ? $signed(regsB_91_re) : $signed(_GEN_7502); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7504 = 8'h1e == _T_24 ? $signed(32'sh0) : $signed(_GEN_7503); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7505 = 8'h1f == _T_24 ? $signed(32'sh0) : $signed(_GEN_7504); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7506 = 8'h20 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7505); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7507 = 8'h21 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7506); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7508 = 8'h22 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7507); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7509 = 8'h23 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7508); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7510 = 8'h24 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7509); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7511 = 8'h25 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7510); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7512 = 8'h26 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7511); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7513 = 8'h27 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7512); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7514 = 8'h28 == _T_24 ? $signed(regsB_2_re) : $signed(_GEN_7513); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7515 = 8'h29 == _T_24 ? $signed(regsB_12_re) : $signed(_GEN_7514); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7516 = 8'h2a == _T_24 ? $signed(regsB_22_re) : $signed(_GEN_7515); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7517 = 8'h2b == _T_24 ? $signed(regsB_32_re) : $signed(_GEN_7516); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7518 = 8'h2c == _T_24 ? $signed(regsB_42_re) : $signed(_GEN_7517); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7519 = 8'h2d == _T_24 ? $signed(regsB_52_re) : $signed(_GEN_7518); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7520 = 8'h2e == _T_24 ? $signed(regsB_62_re) : $signed(_GEN_7519); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7521 = 8'h2f == _T_24 ? $signed(regsB_72_re) : $signed(_GEN_7520); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7522 = 8'h30 == _T_24 ? $signed(regsB_82_re) : $signed(_GEN_7521); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7523 = 8'h31 == _T_24 ? $signed(regsB_92_re) : $signed(_GEN_7522); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7524 = 8'h32 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7523); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7525 = 8'h33 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7524); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7526 = 8'h34 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7525); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7527 = 8'h35 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7526); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7528 = 8'h36 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7527); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7529 = 8'h37 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7528); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7530 = 8'h38 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7529); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7531 = 8'h39 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7530); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7532 = 8'h3a == _T_24 ? $signed(32'sh0) : $signed(_GEN_7531); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7533 = 8'h3b == _T_24 ? $signed(32'sh0) : $signed(_GEN_7532); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7534 = 8'h3c == _T_24 ? $signed(regsB_3_re) : $signed(_GEN_7533); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7535 = 8'h3d == _T_24 ? $signed(regsB_13_re) : $signed(_GEN_7534); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7536 = 8'h3e == _T_24 ? $signed(regsB_23_re) : $signed(_GEN_7535); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7537 = 8'h3f == _T_24 ? $signed(regsB_33_re) : $signed(_GEN_7536); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7538 = 8'h40 == _T_24 ? $signed(regsB_43_re) : $signed(_GEN_7537); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7539 = 8'h41 == _T_24 ? $signed(regsB_53_re) : $signed(_GEN_7538); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7540 = 8'h42 == _T_24 ? $signed(regsB_63_re) : $signed(_GEN_7539); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7541 = 8'h43 == _T_24 ? $signed(regsB_73_re) : $signed(_GEN_7540); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7542 = 8'h44 == _T_24 ? $signed(regsB_83_re) : $signed(_GEN_7541); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7543 = 8'h45 == _T_24 ? $signed(regsB_93_re) : $signed(_GEN_7542); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7544 = 8'h46 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7543); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7545 = 8'h47 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7544); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7546 = 8'h48 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7545); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7547 = 8'h49 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7546); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7548 = 8'h4a == _T_24 ? $signed(32'sh0) : $signed(_GEN_7547); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7549 = 8'h4b == _T_24 ? $signed(32'sh0) : $signed(_GEN_7548); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7550 = 8'h4c == _T_24 ? $signed(32'sh0) : $signed(_GEN_7549); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7551 = 8'h4d == _T_24 ? $signed(32'sh0) : $signed(_GEN_7550); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7552 = 8'h4e == _T_24 ? $signed(32'sh0) : $signed(_GEN_7551); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7553 = 8'h4f == _T_24 ? $signed(32'sh0) : $signed(_GEN_7552); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7554 = 8'h50 == _T_24 ? $signed(regsB_4_re) : $signed(_GEN_7553); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7555 = 8'h51 == _T_24 ? $signed(regsB_14_re) : $signed(_GEN_7554); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7556 = 8'h52 == _T_24 ? $signed(regsB_24_re) : $signed(_GEN_7555); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7557 = 8'h53 == _T_24 ? $signed(regsB_34_re) : $signed(_GEN_7556); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7558 = 8'h54 == _T_24 ? $signed(regsB_44_re) : $signed(_GEN_7557); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7559 = 8'h55 == _T_24 ? $signed(regsB_54_re) : $signed(_GEN_7558); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7560 = 8'h56 == _T_24 ? $signed(regsB_64_re) : $signed(_GEN_7559); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7561 = 8'h57 == _T_24 ? $signed(regsB_74_re) : $signed(_GEN_7560); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7562 = 8'h58 == _T_24 ? $signed(regsB_84_re) : $signed(_GEN_7561); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7563 = 8'h59 == _T_24 ? $signed(regsB_94_re) : $signed(_GEN_7562); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7564 = 8'h5a == _T_24 ? $signed(32'sh0) : $signed(_GEN_7563); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7565 = 8'h5b == _T_24 ? $signed(32'sh0) : $signed(_GEN_7564); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7566 = 8'h5c == _T_24 ? $signed(32'sh0) : $signed(_GEN_7565); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7567 = 8'h5d == _T_24 ? $signed(32'sh0) : $signed(_GEN_7566); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7568 = 8'h5e == _T_24 ? $signed(32'sh0) : $signed(_GEN_7567); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7569 = 8'h5f == _T_24 ? $signed(32'sh0) : $signed(_GEN_7568); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7570 = 8'h60 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7569); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7571 = 8'h61 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7570); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7572 = 8'h62 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7571); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7573 = 8'h63 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7572); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7574 = 8'h64 == _T_24 ? $signed(regsB_5_re) : $signed(_GEN_7573); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7575 = 8'h65 == _T_24 ? $signed(regsB_15_re) : $signed(_GEN_7574); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7576 = 8'h66 == _T_24 ? $signed(regsB_25_re) : $signed(_GEN_7575); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7577 = 8'h67 == _T_24 ? $signed(regsB_35_re) : $signed(_GEN_7576); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7578 = 8'h68 == _T_24 ? $signed(regsB_45_re) : $signed(_GEN_7577); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7579 = 8'h69 == _T_24 ? $signed(regsB_55_re) : $signed(_GEN_7578); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7580 = 8'h6a == _T_24 ? $signed(regsB_65_re) : $signed(_GEN_7579); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7581 = 8'h6b == _T_24 ? $signed(regsB_75_re) : $signed(_GEN_7580); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7582 = 8'h6c == _T_24 ? $signed(regsB_85_re) : $signed(_GEN_7581); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7583 = 8'h6d == _T_24 ? $signed(regsB_95_re) : $signed(_GEN_7582); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7584 = 8'h6e == _T_24 ? $signed(32'sh0) : $signed(_GEN_7583); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7585 = 8'h6f == _T_24 ? $signed(32'sh0) : $signed(_GEN_7584); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7586 = 8'h70 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7585); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7587 = 8'h71 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7586); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7588 = 8'h72 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7587); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7589 = 8'h73 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7588); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7590 = 8'h74 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7589); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7591 = 8'h75 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7590); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7592 = 8'h76 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7591); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7593 = 8'h77 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7592); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7594 = 8'h78 == _T_24 ? $signed(regsB_6_re) : $signed(_GEN_7593); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7595 = 8'h79 == _T_24 ? $signed(regsB_16_re) : $signed(_GEN_7594); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7596 = 8'h7a == _T_24 ? $signed(regsB_26_re) : $signed(_GEN_7595); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7597 = 8'h7b == _T_24 ? $signed(regsB_36_re) : $signed(_GEN_7596); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7598 = 8'h7c == _T_24 ? $signed(regsB_46_re) : $signed(_GEN_7597); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7599 = 8'h7d == _T_24 ? $signed(regsB_56_re) : $signed(_GEN_7598); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7600 = 8'h7e == _T_24 ? $signed(regsB_66_re) : $signed(_GEN_7599); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7601 = 8'h7f == _T_24 ? $signed(regsB_76_re) : $signed(_GEN_7600); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7602 = 8'h80 == _T_24 ? $signed(regsB_86_re) : $signed(_GEN_7601); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7603 = 8'h81 == _T_24 ? $signed(regsB_96_re) : $signed(_GEN_7602); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7604 = 8'h82 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7603); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7605 = 8'h83 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7604); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7606 = 8'h84 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7605); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7607 = 8'h85 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7606); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7608 = 8'h86 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7607); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7609 = 8'h87 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7608); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7610 = 8'h88 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7609); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7611 = 8'h89 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7610); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7612 = 8'h8a == _T_24 ? $signed(32'sh0) : $signed(_GEN_7611); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7613 = 8'h8b == _T_24 ? $signed(32'sh0) : $signed(_GEN_7612); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7614 = 8'h8c == _T_24 ? $signed(regsB_7_re) : $signed(_GEN_7613); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7615 = 8'h8d == _T_24 ? $signed(regsB_17_re) : $signed(_GEN_7614); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7616 = 8'h8e == _T_24 ? $signed(regsB_27_re) : $signed(_GEN_7615); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7617 = 8'h8f == _T_24 ? $signed(regsB_37_re) : $signed(_GEN_7616); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7618 = 8'h90 == _T_24 ? $signed(regsB_47_re) : $signed(_GEN_7617); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7619 = 8'h91 == _T_24 ? $signed(regsB_57_re) : $signed(_GEN_7618); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7620 = 8'h92 == _T_24 ? $signed(regsB_67_re) : $signed(_GEN_7619); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7621 = 8'h93 == _T_24 ? $signed(regsB_77_re) : $signed(_GEN_7620); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7622 = 8'h94 == _T_24 ? $signed(regsB_87_re) : $signed(_GEN_7621); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7623 = 8'h95 == _T_24 ? $signed(regsB_97_re) : $signed(_GEN_7622); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7624 = 8'h96 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7623); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7625 = 8'h97 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7624); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7626 = 8'h98 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7625); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7627 = 8'h99 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7626); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7628 = 8'h9a == _T_24 ? $signed(32'sh0) : $signed(_GEN_7627); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7629 = 8'h9b == _T_24 ? $signed(32'sh0) : $signed(_GEN_7628); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7630 = 8'h9c == _T_24 ? $signed(32'sh0) : $signed(_GEN_7629); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7631 = 8'h9d == _T_24 ? $signed(32'sh0) : $signed(_GEN_7630); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7632 = 8'h9e == _T_24 ? $signed(32'sh0) : $signed(_GEN_7631); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7633 = 8'h9f == _T_24 ? $signed(32'sh0) : $signed(_GEN_7632); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7634 = 8'ha0 == _T_24 ? $signed(regsB_8_re) : $signed(_GEN_7633); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7635 = 8'ha1 == _T_24 ? $signed(regsB_18_re) : $signed(_GEN_7634); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7636 = 8'ha2 == _T_24 ? $signed(regsB_28_re) : $signed(_GEN_7635); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7637 = 8'ha3 == _T_24 ? $signed(regsB_38_re) : $signed(_GEN_7636); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7638 = 8'ha4 == _T_24 ? $signed(regsB_48_re) : $signed(_GEN_7637); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7639 = 8'ha5 == _T_24 ? $signed(regsB_58_re) : $signed(_GEN_7638); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7640 = 8'ha6 == _T_24 ? $signed(regsB_68_re) : $signed(_GEN_7639); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7641 = 8'ha7 == _T_24 ? $signed(regsB_78_re) : $signed(_GEN_7640); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7642 = 8'ha8 == _T_24 ? $signed(regsB_88_re) : $signed(_GEN_7641); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7643 = 8'ha9 == _T_24 ? $signed(regsB_98_re) : $signed(_GEN_7642); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7644 = 8'haa == _T_24 ? $signed(32'sh0) : $signed(_GEN_7643); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7645 = 8'hab == _T_24 ? $signed(32'sh0) : $signed(_GEN_7644); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7646 = 8'hac == _T_24 ? $signed(32'sh0) : $signed(_GEN_7645); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7647 = 8'had == _T_24 ? $signed(32'sh0) : $signed(_GEN_7646); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7648 = 8'hae == _T_24 ? $signed(32'sh0) : $signed(_GEN_7647); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7649 = 8'haf == _T_24 ? $signed(32'sh0) : $signed(_GEN_7648); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7650 = 8'hb0 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7649); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7651 = 8'hb1 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7650); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7652 = 8'hb2 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7651); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7653 = 8'hb3 == _T_24 ? $signed(32'sh0) : $signed(_GEN_7652); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7654 = 8'hb4 == _T_24 ? $signed(regsB_9_re) : $signed(_GEN_7653); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7655 = 8'hb5 == _T_24 ? $signed(regsB_19_re) : $signed(_GEN_7654); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7656 = 8'hb6 == _T_24 ? $signed(regsB_29_re) : $signed(_GEN_7655); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7657 = 8'hb7 == _T_24 ? $signed(regsB_39_re) : $signed(_GEN_7656); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7658 = 8'hb8 == _T_24 ? $signed(regsB_49_re) : $signed(_GEN_7657); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7659 = 8'hb9 == _T_24 ? $signed(regsB_59_re) : $signed(_GEN_7658); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7660 = 8'hba == _T_24 ? $signed(regsB_69_re) : $signed(_GEN_7659); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7661 = 8'hbb == _T_24 ? $signed(regsB_79_re) : $signed(_GEN_7660); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7662 = 8'hbc == _T_24 ? $signed(regsB_89_re) : $signed(_GEN_7661); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7663 = 8'hbd == _T_24 ? $signed(regsB_99_re) : $signed(_GEN_7662); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7665 = 8'h1 == _T_27[7:0] ? $signed(regsB_10_im) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7666 = 8'h2 == _T_27[7:0] ? $signed(regsB_20_im) : $signed(_GEN_7665); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7667 = 8'h3 == _T_27[7:0] ? $signed(regsB_30_im) : $signed(_GEN_7666); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7668 = 8'h4 == _T_27[7:0] ? $signed(regsB_40_im) : $signed(_GEN_7667); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7669 = 8'h5 == _T_27[7:0] ? $signed(regsB_50_im) : $signed(_GEN_7668); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7670 = 8'h6 == _T_27[7:0] ? $signed(regsB_60_im) : $signed(_GEN_7669); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7671 = 8'h7 == _T_27[7:0] ? $signed(regsB_70_im) : $signed(_GEN_7670); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7672 = 8'h8 == _T_27[7:0] ? $signed(regsB_80_im) : $signed(_GEN_7671); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7673 = 8'h9 == _T_27[7:0] ? $signed(regsB_90_im) : $signed(_GEN_7672); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7674 = 8'ha == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7673); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7675 = 8'hb == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7674); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7676 = 8'hc == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7675); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7677 = 8'hd == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7676); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7678 = 8'he == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7677); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7679 = 8'hf == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7678); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7680 = 8'h10 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7679); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7681 = 8'h11 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7680); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7682 = 8'h12 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7681); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7683 = 8'h13 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7682); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7684 = 8'h14 == _T_27[7:0] ? $signed(regsB_1_im) : $signed(_GEN_7683); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7685 = 8'h15 == _T_27[7:0] ? $signed(regsB_11_im) : $signed(_GEN_7684); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7686 = 8'h16 == _T_27[7:0] ? $signed(regsB_21_im) : $signed(_GEN_7685); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7687 = 8'h17 == _T_27[7:0] ? $signed(regsB_31_im) : $signed(_GEN_7686); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7688 = 8'h18 == _T_27[7:0] ? $signed(regsB_41_im) : $signed(_GEN_7687); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7689 = 8'h19 == _T_27[7:0] ? $signed(regsB_51_im) : $signed(_GEN_7688); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7690 = 8'h1a == _T_27[7:0] ? $signed(regsB_61_im) : $signed(_GEN_7689); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7691 = 8'h1b == _T_27[7:0] ? $signed(regsB_71_im) : $signed(_GEN_7690); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7692 = 8'h1c == _T_27[7:0] ? $signed(regsB_81_im) : $signed(_GEN_7691); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7693 = 8'h1d == _T_27[7:0] ? $signed(regsB_91_im) : $signed(_GEN_7692); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7694 = 8'h1e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7693); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7695 = 8'h1f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7694); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7696 = 8'h20 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7695); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7697 = 8'h21 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7696); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7698 = 8'h22 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7697); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7699 = 8'h23 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7698); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7700 = 8'h24 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7699); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7701 = 8'h25 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7700); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7702 = 8'h26 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7701); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7703 = 8'h27 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7702); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7704 = 8'h28 == _T_27[7:0] ? $signed(regsB_2_im) : $signed(_GEN_7703); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7705 = 8'h29 == _T_27[7:0] ? $signed(regsB_12_im) : $signed(_GEN_7704); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7706 = 8'h2a == _T_27[7:0] ? $signed(regsB_22_im) : $signed(_GEN_7705); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7707 = 8'h2b == _T_27[7:0] ? $signed(regsB_32_im) : $signed(_GEN_7706); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7708 = 8'h2c == _T_27[7:0] ? $signed(regsB_42_im) : $signed(_GEN_7707); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7709 = 8'h2d == _T_27[7:0] ? $signed(regsB_52_im) : $signed(_GEN_7708); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7710 = 8'h2e == _T_27[7:0] ? $signed(regsB_62_im) : $signed(_GEN_7709); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7711 = 8'h2f == _T_27[7:0] ? $signed(regsB_72_im) : $signed(_GEN_7710); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7712 = 8'h30 == _T_27[7:0] ? $signed(regsB_82_im) : $signed(_GEN_7711); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7713 = 8'h31 == _T_27[7:0] ? $signed(regsB_92_im) : $signed(_GEN_7712); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7714 = 8'h32 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7713); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7715 = 8'h33 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7714); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7716 = 8'h34 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7715); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7717 = 8'h35 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7716); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7718 = 8'h36 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7717); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7719 = 8'h37 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7718); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7720 = 8'h38 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7719); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7721 = 8'h39 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7720); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7722 = 8'h3a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7721); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7723 = 8'h3b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7722); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7724 = 8'h3c == _T_27[7:0] ? $signed(regsB_3_im) : $signed(_GEN_7723); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7725 = 8'h3d == _T_27[7:0] ? $signed(regsB_13_im) : $signed(_GEN_7724); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7726 = 8'h3e == _T_27[7:0] ? $signed(regsB_23_im) : $signed(_GEN_7725); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7727 = 8'h3f == _T_27[7:0] ? $signed(regsB_33_im) : $signed(_GEN_7726); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7728 = 8'h40 == _T_27[7:0] ? $signed(regsB_43_im) : $signed(_GEN_7727); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7729 = 8'h41 == _T_27[7:0] ? $signed(regsB_53_im) : $signed(_GEN_7728); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7730 = 8'h42 == _T_27[7:0] ? $signed(regsB_63_im) : $signed(_GEN_7729); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7731 = 8'h43 == _T_27[7:0] ? $signed(regsB_73_im) : $signed(_GEN_7730); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7732 = 8'h44 == _T_27[7:0] ? $signed(regsB_83_im) : $signed(_GEN_7731); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7733 = 8'h45 == _T_27[7:0] ? $signed(regsB_93_im) : $signed(_GEN_7732); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7734 = 8'h46 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7733); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7735 = 8'h47 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7734); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7736 = 8'h48 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7735); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7737 = 8'h49 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7736); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7738 = 8'h4a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7737); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7739 = 8'h4b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7738); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7740 = 8'h4c == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7739); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7741 = 8'h4d == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7740); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7742 = 8'h4e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7741); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7743 = 8'h4f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7742); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7744 = 8'h50 == _T_27[7:0] ? $signed(regsB_4_im) : $signed(_GEN_7743); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7745 = 8'h51 == _T_27[7:0] ? $signed(regsB_14_im) : $signed(_GEN_7744); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7746 = 8'h52 == _T_27[7:0] ? $signed(regsB_24_im) : $signed(_GEN_7745); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7747 = 8'h53 == _T_27[7:0] ? $signed(regsB_34_im) : $signed(_GEN_7746); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7748 = 8'h54 == _T_27[7:0] ? $signed(regsB_44_im) : $signed(_GEN_7747); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7749 = 8'h55 == _T_27[7:0] ? $signed(regsB_54_im) : $signed(_GEN_7748); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7750 = 8'h56 == _T_27[7:0] ? $signed(regsB_64_im) : $signed(_GEN_7749); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7751 = 8'h57 == _T_27[7:0] ? $signed(regsB_74_im) : $signed(_GEN_7750); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7752 = 8'h58 == _T_27[7:0] ? $signed(regsB_84_im) : $signed(_GEN_7751); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7753 = 8'h59 == _T_27[7:0] ? $signed(regsB_94_im) : $signed(_GEN_7752); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7754 = 8'h5a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7753); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7755 = 8'h5b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7754); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7756 = 8'h5c == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7755); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7757 = 8'h5d == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7756); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7758 = 8'h5e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7757); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7759 = 8'h5f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7758); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7760 = 8'h60 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7759); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7761 = 8'h61 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7760); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7762 = 8'h62 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7761); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7763 = 8'h63 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7762); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7764 = 8'h64 == _T_27[7:0] ? $signed(regsB_5_im) : $signed(_GEN_7763); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7765 = 8'h65 == _T_27[7:0] ? $signed(regsB_15_im) : $signed(_GEN_7764); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7766 = 8'h66 == _T_27[7:0] ? $signed(regsB_25_im) : $signed(_GEN_7765); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7767 = 8'h67 == _T_27[7:0] ? $signed(regsB_35_im) : $signed(_GEN_7766); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7768 = 8'h68 == _T_27[7:0] ? $signed(regsB_45_im) : $signed(_GEN_7767); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7769 = 8'h69 == _T_27[7:0] ? $signed(regsB_55_im) : $signed(_GEN_7768); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7770 = 8'h6a == _T_27[7:0] ? $signed(regsB_65_im) : $signed(_GEN_7769); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7771 = 8'h6b == _T_27[7:0] ? $signed(regsB_75_im) : $signed(_GEN_7770); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7772 = 8'h6c == _T_27[7:0] ? $signed(regsB_85_im) : $signed(_GEN_7771); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7773 = 8'h6d == _T_27[7:0] ? $signed(regsB_95_im) : $signed(_GEN_7772); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7774 = 8'h6e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7773); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7775 = 8'h6f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7774); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7776 = 8'h70 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7775); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7777 = 8'h71 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7776); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7778 = 8'h72 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7777); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7779 = 8'h73 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7778); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7780 = 8'h74 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7779); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7781 = 8'h75 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7780); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7782 = 8'h76 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7781); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7783 = 8'h77 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7782); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7784 = 8'h78 == _T_27[7:0] ? $signed(regsB_6_im) : $signed(_GEN_7783); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7785 = 8'h79 == _T_27[7:0] ? $signed(regsB_16_im) : $signed(_GEN_7784); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7786 = 8'h7a == _T_27[7:0] ? $signed(regsB_26_im) : $signed(_GEN_7785); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7787 = 8'h7b == _T_27[7:0] ? $signed(regsB_36_im) : $signed(_GEN_7786); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7788 = 8'h7c == _T_27[7:0] ? $signed(regsB_46_im) : $signed(_GEN_7787); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7789 = 8'h7d == _T_27[7:0] ? $signed(regsB_56_im) : $signed(_GEN_7788); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7790 = 8'h7e == _T_27[7:0] ? $signed(regsB_66_im) : $signed(_GEN_7789); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7791 = 8'h7f == _T_27[7:0] ? $signed(regsB_76_im) : $signed(_GEN_7790); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7792 = 8'h80 == _T_27[7:0] ? $signed(regsB_86_im) : $signed(_GEN_7791); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7793 = 8'h81 == _T_27[7:0] ? $signed(regsB_96_im) : $signed(_GEN_7792); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7794 = 8'h82 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7793); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7795 = 8'h83 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7794); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7796 = 8'h84 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7795); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7797 = 8'h85 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7796); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7798 = 8'h86 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7797); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7799 = 8'h87 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7798); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7800 = 8'h88 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7799); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7801 = 8'h89 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7800); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7802 = 8'h8a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7801); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7803 = 8'h8b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7802); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7804 = 8'h8c == _T_27[7:0] ? $signed(regsB_7_im) : $signed(_GEN_7803); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7805 = 8'h8d == _T_27[7:0] ? $signed(regsB_17_im) : $signed(_GEN_7804); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7806 = 8'h8e == _T_27[7:0] ? $signed(regsB_27_im) : $signed(_GEN_7805); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7807 = 8'h8f == _T_27[7:0] ? $signed(regsB_37_im) : $signed(_GEN_7806); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7808 = 8'h90 == _T_27[7:0] ? $signed(regsB_47_im) : $signed(_GEN_7807); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7809 = 8'h91 == _T_27[7:0] ? $signed(regsB_57_im) : $signed(_GEN_7808); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7810 = 8'h92 == _T_27[7:0] ? $signed(regsB_67_im) : $signed(_GEN_7809); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7811 = 8'h93 == _T_27[7:0] ? $signed(regsB_77_im) : $signed(_GEN_7810); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7812 = 8'h94 == _T_27[7:0] ? $signed(regsB_87_im) : $signed(_GEN_7811); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7813 = 8'h95 == _T_27[7:0] ? $signed(regsB_97_im) : $signed(_GEN_7812); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7814 = 8'h96 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7813); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7815 = 8'h97 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7814); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7816 = 8'h98 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7815); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7817 = 8'h99 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7816); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7818 = 8'h9a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7817); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7819 = 8'h9b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7818); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7820 = 8'h9c == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7819); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7821 = 8'h9d == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7820); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7822 = 8'h9e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7821); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7823 = 8'h9f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7822); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7824 = 8'ha0 == _T_27[7:0] ? $signed(regsB_8_im) : $signed(_GEN_7823); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7825 = 8'ha1 == _T_27[7:0] ? $signed(regsB_18_im) : $signed(_GEN_7824); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7826 = 8'ha2 == _T_27[7:0] ? $signed(regsB_28_im) : $signed(_GEN_7825); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7827 = 8'ha3 == _T_27[7:0] ? $signed(regsB_38_im) : $signed(_GEN_7826); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7828 = 8'ha4 == _T_27[7:0] ? $signed(regsB_48_im) : $signed(_GEN_7827); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7829 = 8'ha5 == _T_27[7:0] ? $signed(regsB_58_im) : $signed(_GEN_7828); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7830 = 8'ha6 == _T_27[7:0] ? $signed(regsB_68_im) : $signed(_GEN_7829); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7831 = 8'ha7 == _T_27[7:0] ? $signed(regsB_78_im) : $signed(_GEN_7830); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7832 = 8'ha8 == _T_27[7:0] ? $signed(regsB_88_im) : $signed(_GEN_7831); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7833 = 8'ha9 == _T_27[7:0] ? $signed(regsB_98_im) : $signed(_GEN_7832); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7834 = 8'haa == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7833); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7835 = 8'hab == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7834); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7836 = 8'hac == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7835); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7837 = 8'had == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7836); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7838 = 8'hae == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7837); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7839 = 8'haf == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7838); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7840 = 8'hb0 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7839); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7841 = 8'hb1 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7840); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7842 = 8'hb2 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7841); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7843 = 8'hb3 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7842); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7844 = 8'hb4 == _T_27[7:0] ? $signed(regsB_9_im) : $signed(_GEN_7843); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7845 = 8'hb5 == _T_27[7:0] ? $signed(regsB_19_im) : $signed(_GEN_7844); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7846 = 8'hb6 == _T_27[7:0] ? $signed(regsB_29_im) : $signed(_GEN_7845); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7847 = 8'hb7 == _T_27[7:0] ? $signed(regsB_39_im) : $signed(_GEN_7846); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7848 = 8'hb8 == _T_27[7:0] ? $signed(regsB_49_im) : $signed(_GEN_7847); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7849 = 8'hb9 == _T_27[7:0] ? $signed(regsB_59_im) : $signed(_GEN_7848); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7850 = 8'hba == _T_27[7:0] ? $signed(regsB_69_im) : $signed(_GEN_7849); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7851 = 8'hbb == _T_27[7:0] ? $signed(regsB_79_im) : $signed(_GEN_7850); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7852 = 8'hbc == _T_27[7:0] ? $signed(regsB_89_im) : $signed(_GEN_7851); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7853 = 8'hbd == _T_27[7:0] ? $signed(regsB_99_im) : $signed(_GEN_7852); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7855 = 8'h1 == _T_27[7:0] ? $signed(regsB_10_re) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7856 = 8'h2 == _T_27[7:0] ? $signed(regsB_20_re) : $signed(_GEN_7855); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7857 = 8'h3 == _T_27[7:0] ? $signed(regsB_30_re) : $signed(_GEN_7856); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7858 = 8'h4 == _T_27[7:0] ? $signed(regsB_40_re) : $signed(_GEN_7857); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7859 = 8'h5 == _T_27[7:0] ? $signed(regsB_50_re) : $signed(_GEN_7858); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7860 = 8'h6 == _T_27[7:0] ? $signed(regsB_60_re) : $signed(_GEN_7859); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7861 = 8'h7 == _T_27[7:0] ? $signed(regsB_70_re) : $signed(_GEN_7860); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7862 = 8'h8 == _T_27[7:0] ? $signed(regsB_80_re) : $signed(_GEN_7861); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7863 = 8'h9 == _T_27[7:0] ? $signed(regsB_90_re) : $signed(_GEN_7862); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7864 = 8'ha == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7863); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7865 = 8'hb == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7864); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7866 = 8'hc == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7865); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7867 = 8'hd == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7866); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7868 = 8'he == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7867); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7869 = 8'hf == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7868); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7870 = 8'h10 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7869); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7871 = 8'h11 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7870); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7872 = 8'h12 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7871); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7873 = 8'h13 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7872); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7874 = 8'h14 == _T_27[7:0] ? $signed(regsB_1_re) : $signed(_GEN_7873); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7875 = 8'h15 == _T_27[7:0] ? $signed(regsB_11_re) : $signed(_GEN_7874); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7876 = 8'h16 == _T_27[7:0] ? $signed(regsB_21_re) : $signed(_GEN_7875); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7877 = 8'h17 == _T_27[7:0] ? $signed(regsB_31_re) : $signed(_GEN_7876); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7878 = 8'h18 == _T_27[7:0] ? $signed(regsB_41_re) : $signed(_GEN_7877); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7879 = 8'h19 == _T_27[7:0] ? $signed(regsB_51_re) : $signed(_GEN_7878); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7880 = 8'h1a == _T_27[7:0] ? $signed(regsB_61_re) : $signed(_GEN_7879); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7881 = 8'h1b == _T_27[7:0] ? $signed(regsB_71_re) : $signed(_GEN_7880); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7882 = 8'h1c == _T_27[7:0] ? $signed(regsB_81_re) : $signed(_GEN_7881); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7883 = 8'h1d == _T_27[7:0] ? $signed(regsB_91_re) : $signed(_GEN_7882); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7884 = 8'h1e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7883); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7885 = 8'h1f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7884); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7886 = 8'h20 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7885); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7887 = 8'h21 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7886); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7888 = 8'h22 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7887); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7889 = 8'h23 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7888); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7890 = 8'h24 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7889); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7891 = 8'h25 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7890); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7892 = 8'h26 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7891); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7893 = 8'h27 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7892); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7894 = 8'h28 == _T_27[7:0] ? $signed(regsB_2_re) : $signed(_GEN_7893); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7895 = 8'h29 == _T_27[7:0] ? $signed(regsB_12_re) : $signed(_GEN_7894); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7896 = 8'h2a == _T_27[7:0] ? $signed(regsB_22_re) : $signed(_GEN_7895); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7897 = 8'h2b == _T_27[7:0] ? $signed(regsB_32_re) : $signed(_GEN_7896); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7898 = 8'h2c == _T_27[7:0] ? $signed(regsB_42_re) : $signed(_GEN_7897); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7899 = 8'h2d == _T_27[7:0] ? $signed(regsB_52_re) : $signed(_GEN_7898); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7900 = 8'h2e == _T_27[7:0] ? $signed(regsB_62_re) : $signed(_GEN_7899); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7901 = 8'h2f == _T_27[7:0] ? $signed(regsB_72_re) : $signed(_GEN_7900); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7902 = 8'h30 == _T_27[7:0] ? $signed(regsB_82_re) : $signed(_GEN_7901); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7903 = 8'h31 == _T_27[7:0] ? $signed(regsB_92_re) : $signed(_GEN_7902); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7904 = 8'h32 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7903); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7905 = 8'h33 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7904); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7906 = 8'h34 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7905); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7907 = 8'h35 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7906); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7908 = 8'h36 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7907); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7909 = 8'h37 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7908); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7910 = 8'h38 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7909); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7911 = 8'h39 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7910); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7912 = 8'h3a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7911); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7913 = 8'h3b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7912); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7914 = 8'h3c == _T_27[7:0] ? $signed(regsB_3_re) : $signed(_GEN_7913); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7915 = 8'h3d == _T_27[7:0] ? $signed(regsB_13_re) : $signed(_GEN_7914); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7916 = 8'h3e == _T_27[7:0] ? $signed(regsB_23_re) : $signed(_GEN_7915); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7917 = 8'h3f == _T_27[7:0] ? $signed(regsB_33_re) : $signed(_GEN_7916); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7918 = 8'h40 == _T_27[7:0] ? $signed(regsB_43_re) : $signed(_GEN_7917); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7919 = 8'h41 == _T_27[7:0] ? $signed(regsB_53_re) : $signed(_GEN_7918); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7920 = 8'h42 == _T_27[7:0] ? $signed(regsB_63_re) : $signed(_GEN_7919); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7921 = 8'h43 == _T_27[7:0] ? $signed(regsB_73_re) : $signed(_GEN_7920); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7922 = 8'h44 == _T_27[7:0] ? $signed(regsB_83_re) : $signed(_GEN_7921); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7923 = 8'h45 == _T_27[7:0] ? $signed(regsB_93_re) : $signed(_GEN_7922); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7924 = 8'h46 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7923); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7925 = 8'h47 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7924); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7926 = 8'h48 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7925); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7927 = 8'h49 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7926); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7928 = 8'h4a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7927); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7929 = 8'h4b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7928); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7930 = 8'h4c == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7929); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7931 = 8'h4d == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7930); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7932 = 8'h4e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7931); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7933 = 8'h4f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7932); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7934 = 8'h50 == _T_27[7:0] ? $signed(regsB_4_re) : $signed(_GEN_7933); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7935 = 8'h51 == _T_27[7:0] ? $signed(regsB_14_re) : $signed(_GEN_7934); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7936 = 8'h52 == _T_27[7:0] ? $signed(regsB_24_re) : $signed(_GEN_7935); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7937 = 8'h53 == _T_27[7:0] ? $signed(regsB_34_re) : $signed(_GEN_7936); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7938 = 8'h54 == _T_27[7:0] ? $signed(regsB_44_re) : $signed(_GEN_7937); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7939 = 8'h55 == _T_27[7:0] ? $signed(regsB_54_re) : $signed(_GEN_7938); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7940 = 8'h56 == _T_27[7:0] ? $signed(regsB_64_re) : $signed(_GEN_7939); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7941 = 8'h57 == _T_27[7:0] ? $signed(regsB_74_re) : $signed(_GEN_7940); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7942 = 8'h58 == _T_27[7:0] ? $signed(regsB_84_re) : $signed(_GEN_7941); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7943 = 8'h59 == _T_27[7:0] ? $signed(regsB_94_re) : $signed(_GEN_7942); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7944 = 8'h5a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7943); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7945 = 8'h5b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7944); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7946 = 8'h5c == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7945); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7947 = 8'h5d == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7946); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7948 = 8'h5e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7947); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7949 = 8'h5f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7948); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7950 = 8'h60 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7949); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7951 = 8'h61 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7950); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7952 = 8'h62 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7951); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7953 = 8'h63 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7952); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7954 = 8'h64 == _T_27[7:0] ? $signed(regsB_5_re) : $signed(_GEN_7953); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7955 = 8'h65 == _T_27[7:0] ? $signed(regsB_15_re) : $signed(_GEN_7954); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7956 = 8'h66 == _T_27[7:0] ? $signed(regsB_25_re) : $signed(_GEN_7955); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7957 = 8'h67 == _T_27[7:0] ? $signed(regsB_35_re) : $signed(_GEN_7956); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7958 = 8'h68 == _T_27[7:0] ? $signed(regsB_45_re) : $signed(_GEN_7957); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7959 = 8'h69 == _T_27[7:0] ? $signed(regsB_55_re) : $signed(_GEN_7958); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7960 = 8'h6a == _T_27[7:0] ? $signed(regsB_65_re) : $signed(_GEN_7959); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7961 = 8'h6b == _T_27[7:0] ? $signed(regsB_75_re) : $signed(_GEN_7960); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7962 = 8'h6c == _T_27[7:0] ? $signed(regsB_85_re) : $signed(_GEN_7961); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7963 = 8'h6d == _T_27[7:0] ? $signed(regsB_95_re) : $signed(_GEN_7962); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7964 = 8'h6e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7963); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7965 = 8'h6f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7964); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7966 = 8'h70 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7965); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7967 = 8'h71 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7966); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7968 = 8'h72 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7967); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7969 = 8'h73 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7968); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7970 = 8'h74 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7969); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7971 = 8'h75 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7970); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7972 = 8'h76 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7971); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7973 = 8'h77 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7972); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7974 = 8'h78 == _T_27[7:0] ? $signed(regsB_6_re) : $signed(_GEN_7973); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7975 = 8'h79 == _T_27[7:0] ? $signed(regsB_16_re) : $signed(_GEN_7974); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7976 = 8'h7a == _T_27[7:0] ? $signed(regsB_26_re) : $signed(_GEN_7975); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7977 = 8'h7b == _T_27[7:0] ? $signed(regsB_36_re) : $signed(_GEN_7976); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7978 = 8'h7c == _T_27[7:0] ? $signed(regsB_46_re) : $signed(_GEN_7977); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7979 = 8'h7d == _T_27[7:0] ? $signed(regsB_56_re) : $signed(_GEN_7978); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7980 = 8'h7e == _T_27[7:0] ? $signed(regsB_66_re) : $signed(_GEN_7979); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7981 = 8'h7f == _T_27[7:0] ? $signed(regsB_76_re) : $signed(_GEN_7980); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7982 = 8'h80 == _T_27[7:0] ? $signed(regsB_86_re) : $signed(_GEN_7981); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7983 = 8'h81 == _T_27[7:0] ? $signed(regsB_96_re) : $signed(_GEN_7982); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7984 = 8'h82 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7983); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7985 = 8'h83 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7984); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7986 = 8'h84 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7985); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7987 = 8'h85 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7986); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7988 = 8'h86 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7987); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7989 = 8'h87 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7988); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7990 = 8'h88 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7989); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7991 = 8'h89 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7990); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7992 = 8'h8a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7991); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7993 = 8'h8b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_7992); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7994 = 8'h8c == _T_27[7:0] ? $signed(regsB_7_re) : $signed(_GEN_7993); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7995 = 8'h8d == _T_27[7:0] ? $signed(regsB_17_re) : $signed(_GEN_7994); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7996 = 8'h8e == _T_27[7:0] ? $signed(regsB_27_re) : $signed(_GEN_7995); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7997 = 8'h8f == _T_27[7:0] ? $signed(regsB_37_re) : $signed(_GEN_7996); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7998 = 8'h90 == _T_27[7:0] ? $signed(regsB_47_re) : $signed(_GEN_7997); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_7999 = 8'h91 == _T_27[7:0] ? $signed(regsB_57_re) : $signed(_GEN_7998); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8000 = 8'h92 == _T_27[7:0] ? $signed(regsB_67_re) : $signed(_GEN_7999); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8001 = 8'h93 == _T_27[7:0] ? $signed(regsB_77_re) : $signed(_GEN_8000); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8002 = 8'h94 == _T_27[7:0] ? $signed(regsB_87_re) : $signed(_GEN_8001); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8003 = 8'h95 == _T_27[7:0] ? $signed(regsB_97_re) : $signed(_GEN_8002); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8004 = 8'h96 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8003); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8005 = 8'h97 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8004); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8006 = 8'h98 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8005); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8007 = 8'h99 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8006); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8008 = 8'h9a == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8007); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8009 = 8'h9b == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8008); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8010 = 8'h9c == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8009); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8011 = 8'h9d == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8010); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8012 = 8'h9e == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8011); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8013 = 8'h9f == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8012); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8014 = 8'ha0 == _T_27[7:0] ? $signed(regsB_8_re) : $signed(_GEN_8013); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8015 = 8'ha1 == _T_27[7:0] ? $signed(regsB_18_re) : $signed(_GEN_8014); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8016 = 8'ha2 == _T_27[7:0] ? $signed(regsB_28_re) : $signed(_GEN_8015); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8017 = 8'ha3 == _T_27[7:0] ? $signed(regsB_38_re) : $signed(_GEN_8016); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8018 = 8'ha4 == _T_27[7:0] ? $signed(regsB_48_re) : $signed(_GEN_8017); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8019 = 8'ha5 == _T_27[7:0] ? $signed(regsB_58_re) : $signed(_GEN_8018); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8020 = 8'ha6 == _T_27[7:0] ? $signed(regsB_68_re) : $signed(_GEN_8019); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8021 = 8'ha7 == _T_27[7:0] ? $signed(regsB_78_re) : $signed(_GEN_8020); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8022 = 8'ha8 == _T_27[7:0] ? $signed(regsB_88_re) : $signed(_GEN_8021); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8023 = 8'ha9 == _T_27[7:0] ? $signed(regsB_98_re) : $signed(_GEN_8022); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8024 = 8'haa == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8023); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8025 = 8'hab == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8024); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8026 = 8'hac == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8025); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8027 = 8'had == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8026); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8028 = 8'hae == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8027); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8029 = 8'haf == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8028); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8030 = 8'hb0 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8029); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8031 = 8'hb1 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8030); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8032 = 8'hb2 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8031); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8033 = 8'hb3 == _T_27[7:0] ? $signed(32'sh0) : $signed(_GEN_8032); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8034 = 8'hb4 == _T_27[7:0] ? $signed(regsB_9_re) : $signed(_GEN_8033); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8035 = 8'hb5 == _T_27[7:0] ? $signed(regsB_19_re) : $signed(_GEN_8034); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8036 = 8'hb6 == _T_27[7:0] ? $signed(regsB_29_re) : $signed(_GEN_8035); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8037 = 8'hb7 == _T_27[7:0] ? $signed(regsB_39_re) : $signed(_GEN_8036); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8038 = 8'hb8 == _T_27[7:0] ? $signed(regsB_49_re) : $signed(_GEN_8037); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8039 = 8'hb9 == _T_27[7:0] ? $signed(regsB_59_re) : $signed(_GEN_8038); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8040 = 8'hba == _T_27[7:0] ? $signed(regsB_69_re) : $signed(_GEN_8039); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8041 = 8'hbb == _T_27[7:0] ? $signed(regsB_79_re) : $signed(_GEN_8040); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8042 = 8'hbc == _T_27[7:0] ? $signed(regsB_89_re) : $signed(_GEN_8041); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8043 = 8'hbd == _T_27[7:0] ? $signed(regsB_99_re) : $signed(_GEN_8042); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8045 = 8'h1 == _T_31[7:0] ? $signed(regsB_10_im) : $signed(regsB_0_im); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8046 = 8'h2 == _T_31[7:0] ? $signed(regsB_20_im) : $signed(_GEN_8045); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8047 = 8'h3 == _T_31[7:0] ? $signed(regsB_30_im) : $signed(_GEN_8046); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8048 = 8'h4 == _T_31[7:0] ? $signed(regsB_40_im) : $signed(_GEN_8047); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8049 = 8'h5 == _T_31[7:0] ? $signed(regsB_50_im) : $signed(_GEN_8048); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8050 = 8'h6 == _T_31[7:0] ? $signed(regsB_60_im) : $signed(_GEN_8049); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8051 = 8'h7 == _T_31[7:0] ? $signed(regsB_70_im) : $signed(_GEN_8050); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8052 = 8'h8 == _T_31[7:0] ? $signed(regsB_80_im) : $signed(_GEN_8051); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8053 = 8'h9 == _T_31[7:0] ? $signed(regsB_90_im) : $signed(_GEN_8052); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8054 = 8'ha == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8053); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8055 = 8'hb == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8054); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8056 = 8'hc == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8055); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8057 = 8'hd == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8056); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8058 = 8'he == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8057); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8059 = 8'hf == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8058); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8060 = 8'h10 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8059); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8061 = 8'h11 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8060); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8062 = 8'h12 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8061); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8063 = 8'h13 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8062); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8064 = 8'h14 == _T_31[7:0] ? $signed(regsB_1_im) : $signed(_GEN_8063); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8065 = 8'h15 == _T_31[7:0] ? $signed(regsB_11_im) : $signed(_GEN_8064); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8066 = 8'h16 == _T_31[7:0] ? $signed(regsB_21_im) : $signed(_GEN_8065); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8067 = 8'h17 == _T_31[7:0] ? $signed(regsB_31_im) : $signed(_GEN_8066); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8068 = 8'h18 == _T_31[7:0] ? $signed(regsB_41_im) : $signed(_GEN_8067); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8069 = 8'h19 == _T_31[7:0] ? $signed(regsB_51_im) : $signed(_GEN_8068); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8070 = 8'h1a == _T_31[7:0] ? $signed(regsB_61_im) : $signed(_GEN_8069); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8071 = 8'h1b == _T_31[7:0] ? $signed(regsB_71_im) : $signed(_GEN_8070); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8072 = 8'h1c == _T_31[7:0] ? $signed(regsB_81_im) : $signed(_GEN_8071); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8073 = 8'h1d == _T_31[7:0] ? $signed(regsB_91_im) : $signed(_GEN_8072); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8074 = 8'h1e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8073); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8075 = 8'h1f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8074); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8076 = 8'h20 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8075); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8077 = 8'h21 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8076); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8078 = 8'h22 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8077); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8079 = 8'h23 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8078); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8080 = 8'h24 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8079); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8081 = 8'h25 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8080); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8082 = 8'h26 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8081); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8083 = 8'h27 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8082); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8084 = 8'h28 == _T_31[7:0] ? $signed(regsB_2_im) : $signed(_GEN_8083); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8085 = 8'h29 == _T_31[7:0] ? $signed(regsB_12_im) : $signed(_GEN_8084); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8086 = 8'h2a == _T_31[7:0] ? $signed(regsB_22_im) : $signed(_GEN_8085); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8087 = 8'h2b == _T_31[7:0] ? $signed(regsB_32_im) : $signed(_GEN_8086); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8088 = 8'h2c == _T_31[7:0] ? $signed(regsB_42_im) : $signed(_GEN_8087); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8089 = 8'h2d == _T_31[7:0] ? $signed(regsB_52_im) : $signed(_GEN_8088); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8090 = 8'h2e == _T_31[7:0] ? $signed(regsB_62_im) : $signed(_GEN_8089); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8091 = 8'h2f == _T_31[7:0] ? $signed(regsB_72_im) : $signed(_GEN_8090); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8092 = 8'h30 == _T_31[7:0] ? $signed(regsB_82_im) : $signed(_GEN_8091); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8093 = 8'h31 == _T_31[7:0] ? $signed(regsB_92_im) : $signed(_GEN_8092); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8094 = 8'h32 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8093); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8095 = 8'h33 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8094); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8096 = 8'h34 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8095); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8097 = 8'h35 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8096); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8098 = 8'h36 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8097); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8099 = 8'h37 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8098); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8100 = 8'h38 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8099); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8101 = 8'h39 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8100); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8102 = 8'h3a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8101); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8103 = 8'h3b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8102); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8104 = 8'h3c == _T_31[7:0] ? $signed(regsB_3_im) : $signed(_GEN_8103); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8105 = 8'h3d == _T_31[7:0] ? $signed(regsB_13_im) : $signed(_GEN_8104); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8106 = 8'h3e == _T_31[7:0] ? $signed(regsB_23_im) : $signed(_GEN_8105); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8107 = 8'h3f == _T_31[7:0] ? $signed(regsB_33_im) : $signed(_GEN_8106); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8108 = 8'h40 == _T_31[7:0] ? $signed(regsB_43_im) : $signed(_GEN_8107); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8109 = 8'h41 == _T_31[7:0] ? $signed(regsB_53_im) : $signed(_GEN_8108); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8110 = 8'h42 == _T_31[7:0] ? $signed(regsB_63_im) : $signed(_GEN_8109); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8111 = 8'h43 == _T_31[7:0] ? $signed(regsB_73_im) : $signed(_GEN_8110); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8112 = 8'h44 == _T_31[7:0] ? $signed(regsB_83_im) : $signed(_GEN_8111); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8113 = 8'h45 == _T_31[7:0] ? $signed(regsB_93_im) : $signed(_GEN_8112); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8114 = 8'h46 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8113); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8115 = 8'h47 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8114); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8116 = 8'h48 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8115); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8117 = 8'h49 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8116); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8118 = 8'h4a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8117); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8119 = 8'h4b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8118); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8120 = 8'h4c == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8119); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8121 = 8'h4d == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8120); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8122 = 8'h4e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8121); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8123 = 8'h4f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8122); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8124 = 8'h50 == _T_31[7:0] ? $signed(regsB_4_im) : $signed(_GEN_8123); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8125 = 8'h51 == _T_31[7:0] ? $signed(regsB_14_im) : $signed(_GEN_8124); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8126 = 8'h52 == _T_31[7:0] ? $signed(regsB_24_im) : $signed(_GEN_8125); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8127 = 8'h53 == _T_31[7:0] ? $signed(regsB_34_im) : $signed(_GEN_8126); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8128 = 8'h54 == _T_31[7:0] ? $signed(regsB_44_im) : $signed(_GEN_8127); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8129 = 8'h55 == _T_31[7:0] ? $signed(regsB_54_im) : $signed(_GEN_8128); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8130 = 8'h56 == _T_31[7:0] ? $signed(regsB_64_im) : $signed(_GEN_8129); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8131 = 8'h57 == _T_31[7:0] ? $signed(regsB_74_im) : $signed(_GEN_8130); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8132 = 8'h58 == _T_31[7:0] ? $signed(regsB_84_im) : $signed(_GEN_8131); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8133 = 8'h59 == _T_31[7:0] ? $signed(regsB_94_im) : $signed(_GEN_8132); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8134 = 8'h5a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8133); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8135 = 8'h5b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8134); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8136 = 8'h5c == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8135); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8137 = 8'h5d == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8136); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8138 = 8'h5e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8137); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8139 = 8'h5f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8138); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8140 = 8'h60 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8139); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8141 = 8'h61 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8140); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8142 = 8'h62 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8141); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8143 = 8'h63 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8142); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8144 = 8'h64 == _T_31[7:0] ? $signed(regsB_5_im) : $signed(_GEN_8143); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8145 = 8'h65 == _T_31[7:0] ? $signed(regsB_15_im) : $signed(_GEN_8144); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8146 = 8'h66 == _T_31[7:0] ? $signed(regsB_25_im) : $signed(_GEN_8145); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8147 = 8'h67 == _T_31[7:0] ? $signed(regsB_35_im) : $signed(_GEN_8146); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8148 = 8'h68 == _T_31[7:0] ? $signed(regsB_45_im) : $signed(_GEN_8147); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8149 = 8'h69 == _T_31[7:0] ? $signed(regsB_55_im) : $signed(_GEN_8148); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8150 = 8'h6a == _T_31[7:0] ? $signed(regsB_65_im) : $signed(_GEN_8149); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8151 = 8'h6b == _T_31[7:0] ? $signed(regsB_75_im) : $signed(_GEN_8150); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8152 = 8'h6c == _T_31[7:0] ? $signed(regsB_85_im) : $signed(_GEN_8151); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8153 = 8'h6d == _T_31[7:0] ? $signed(regsB_95_im) : $signed(_GEN_8152); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8154 = 8'h6e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8153); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8155 = 8'h6f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8154); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8156 = 8'h70 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8155); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8157 = 8'h71 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8156); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8158 = 8'h72 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8157); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8159 = 8'h73 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8158); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8160 = 8'h74 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8159); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8161 = 8'h75 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8160); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8162 = 8'h76 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8161); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8163 = 8'h77 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8162); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8164 = 8'h78 == _T_31[7:0] ? $signed(regsB_6_im) : $signed(_GEN_8163); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8165 = 8'h79 == _T_31[7:0] ? $signed(regsB_16_im) : $signed(_GEN_8164); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8166 = 8'h7a == _T_31[7:0] ? $signed(regsB_26_im) : $signed(_GEN_8165); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8167 = 8'h7b == _T_31[7:0] ? $signed(regsB_36_im) : $signed(_GEN_8166); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8168 = 8'h7c == _T_31[7:0] ? $signed(regsB_46_im) : $signed(_GEN_8167); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8169 = 8'h7d == _T_31[7:0] ? $signed(regsB_56_im) : $signed(_GEN_8168); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8170 = 8'h7e == _T_31[7:0] ? $signed(regsB_66_im) : $signed(_GEN_8169); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8171 = 8'h7f == _T_31[7:0] ? $signed(regsB_76_im) : $signed(_GEN_8170); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8172 = 8'h80 == _T_31[7:0] ? $signed(regsB_86_im) : $signed(_GEN_8171); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8173 = 8'h81 == _T_31[7:0] ? $signed(regsB_96_im) : $signed(_GEN_8172); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8174 = 8'h82 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8173); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8175 = 8'h83 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8174); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8176 = 8'h84 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8175); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8177 = 8'h85 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8176); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8178 = 8'h86 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8177); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8179 = 8'h87 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8178); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8180 = 8'h88 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8179); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8181 = 8'h89 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8180); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8182 = 8'h8a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8181); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8183 = 8'h8b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8182); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8184 = 8'h8c == _T_31[7:0] ? $signed(regsB_7_im) : $signed(_GEN_8183); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8185 = 8'h8d == _T_31[7:0] ? $signed(regsB_17_im) : $signed(_GEN_8184); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8186 = 8'h8e == _T_31[7:0] ? $signed(regsB_27_im) : $signed(_GEN_8185); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8187 = 8'h8f == _T_31[7:0] ? $signed(regsB_37_im) : $signed(_GEN_8186); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8188 = 8'h90 == _T_31[7:0] ? $signed(regsB_47_im) : $signed(_GEN_8187); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8189 = 8'h91 == _T_31[7:0] ? $signed(regsB_57_im) : $signed(_GEN_8188); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8190 = 8'h92 == _T_31[7:0] ? $signed(regsB_67_im) : $signed(_GEN_8189); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8191 = 8'h93 == _T_31[7:0] ? $signed(regsB_77_im) : $signed(_GEN_8190); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8192 = 8'h94 == _T_31[7:0] ? $signed(regsB_87_im) : $signed(_GEN_8191); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8193 = 8'h95 == _T_31[7:0] ? $signed(regsB_97_im) : $signed(_GEN_8192); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8194 = 8'h96 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8193); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8195 = 8'h97 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8194); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8196 = 8'h98 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8195); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8197 = 8'h99 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8196); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8198 = 8'h9a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8197); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8199 = 8'h9b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8198); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8200 = 8'h9c == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8199); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8201 = 8'h9d == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8200); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8202 = 8'h9e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8201); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8203 = 8'h9f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8202); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8204 = 8'ha0 == _T_31[7:0] ? $signed(regsB_8_im) : $signed(_GEN_8203); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8205 = 8'ha1 == _T_31[7:0] ? $signed(regsB_18_im) : $signed(_GEN_8204); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8206 = 8'ha2 == _T_31[7:0] ? $signed(regsB_28_im) : $signed(_GEN_8205); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8207 = 8'ha3 == _T_31[7:0] ? $signed(regsB_38_im) : $signed(_GEN_8206); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8208 = 8'ha4 == _T_31[7:0] ? $signed(regsB_48_im) : $signed(_GEN_8207); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8209 = 8'ha5 == _T_31[7:0] ? $signed(regsB_58_im) : $signed(_GEN_8208); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8210 = 8'ha6 == _T_31[7:0] ? $signed(regsB_68_im) : $signed(_GEN_8209); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8211 = 8'ha7 == _T_31[7:0] ? $signed(regsB_78_im) : $signed(_GEN_8210); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8212 = 8'ha8 == _T_31[7:0] ? $signed(regsB_88_im) : $signed(_GEN_8211); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8213 = 8'ha9 == _T_31[7:0] ? $signed(regsB_98_im) : $signed(_GEN_8212); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8214 = 8'haa == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8213); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8215 = 8'hab == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8214); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8216 = 8'hac == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8215); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8217 = 8'had == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8216); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8218 = 8'hae == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8217); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8219 = 8'haf == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8218); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8220 = 8'hb0 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8219); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8221 = 8'hb1 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8220); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8222 = 8'hb2 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8221); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8223 = 8'hb3 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8222); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8224 = 8'hb4 == _T_31[7:0] ? $signed(regsB_9_im) : $signed(_GEN_8223); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8225 = 8'hb5 == _T_31[7:0] ? $signed(regsB_19_im) : $signed(_GEN_8224); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8226 = 8'hb6 == _T_31[7:0] ? $signed(regsB_29_im) : $signed(_GEN_8225); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8227 = 8'hb7 == _T_31[7:0] ? $signed(regsB_39_im) : $signed(_GEN_8226); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8228 = 8'hb8 == _T_31[7:0] ? $signed(regsB_49_im) : $signed(_GEN_8227); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8229 = 8'hb9 == _T_31[7:0] ? $signed(regsB_59_im) : $signed(_GEN_8228); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8230 = 8'hba == _T_31[7:0] ? $signed(regsB_69_im) : $signed(_GEN_8229); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8231 = 8'hbb == _T_31[7:0] ? $signed(regsB_79_im) : $signed(_GEN_8230); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8232 = 8'hbc == _T_31[7:0] ? $signed(regsB_89_im) : $signed(_GEN_8231); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8233 = 8'hbd == _T_31[7:0] ? $signed(regsB_99_im) : $signed(_GEN_8232); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8235 = 8'h1 == _T_31[7:0] ? $signed(regsB_10_re) : $signed(regsB_0_re); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8236 = 8'h2 == _T_31[7:0] ? $signed(regsB_20_re) : $signed(_GEN_8235); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8237 = 8'h3 == _T_31[7:0] ? $signed(regsB_30_re) : $signed(_GEN_8236); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8238 = 8'h4 == _T_31[7:0] ? $signed(regsB_40_re) : $signed(_GEN_8237); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8239 = 8'h5 == _T_31[7:0] ? $signed(regsB_50_re) : $signed(_GEN_8238); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8240 = 8'h6 == _T_31[7:0] ? $signed(regsB_60_re) : $signed(_GEN_8239); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8241 = 8'h7 == _T_31[7:0] ? $signed(regsB_70_re) : $signed(_GEN_8240); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8242 = 8'h8 == _T_31[7:0] ? $signed(regsB_80_re) : $signed(_GEN_8241); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8243 = 8'h9 == _T_31[7:0] ? $signed(regsB_90_re) : $signed(_GEN_8242); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8244 = 8'ha == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8243); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8245 = 8'hb == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8244); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8246 = 8'hc == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8245); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8247 = 8'hd == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8246); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8248 = 8'he == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8247); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8249 = 8'hf == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8248); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8250 = 8'h10 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8249); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8251 = 8'h11 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8250); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8252 = 8'h12 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8251); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8253 = 8'h13 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8252); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8254 = 8'h14 == _T_31[7:0] ? $signed(regsB_1_re) : $signed(_GEN_8253); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8255 = 8'h15 == _T_31[7:0] ? $signed(regsB_11_re) : $signed(_GEN_8254); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8256 = 8'h16 == _T_31[7:0] ? $signed(regsB_21_re) : $signed(_GEN_8255); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8257 = 8'h17 == _T_31[7:0] ? $signed(regsB_31_re) : $signed(_GEN_8256); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8258 = 8'h18 == _T_31[7:0] ? $signed(regsB_41_re) : $signed(_GEN_8257); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8259 = 8'h19 == _T_31[7:0] ? $signed(regsB_51_re) : $signed(_GEN_8258); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8260 = 8'h1a == _T_31[7:0] ? $signed(regsB_61_re) : $signed(_GEN_8259); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8261 = 8'h1b == _T_31[7:0] ? $signed(regsB_71_re) : $signed(_GEN_8260); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8262 = 8'h1c == _T_31[7:0] ? $signed(regsB_81_re) : $signed(_GEN_8261); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8263 = 8'h1d == _T_31[7:0] ? $signed(regsB_91_re) : $signed(_GEN_8262); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8264 = 8'h1e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8263); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8265 = 8'h1f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8264); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8266 = 8'h20 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8265); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8267 = 8'h21 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8266); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8268 = 8'h22 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8267); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8269 = 8'h23 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8268); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8270 = 8'h24 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8269); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8271 = 8'h25 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8270); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8272 = 8'h26 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8271); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8273 = 8'h27 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8272); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8274 = 8'h28 == _T_31[7:0] ? $signed(regsB_2_re) : $signed(_GEN_8273); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8275 = 8'h29 == _T_31[7:0] ? $signed(regsB_12_re) : $signed(_GEN_8274); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8276 = 8'h2a == _T_31[7:0] ? $signed(regsB_22_re) : $signed(_GEN_8275); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8277 = 8'h2b == _T_31[7:0] ? $signed(regsB_32_re) : $signed(_GEN_8276); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8278 = 8'h2c == _T_31[7:0] ? $signed(regsB_42_re) : $signed(_GEN_8277); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8279 = 8'h2d == _T_31[7:0] ? $signed(regsB_52_re) : $signed(_GEN_8278); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8280 = 8'h2e == _T_31[7:0] ? $signed(regsB_62_re) : $signed(_GEN_8279); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8281 = 8'h2f == _T_31[7:0] ? $signed(regsB_72_re) : $signed(_GEN_8280); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8282 = 8'h30 == _T_31[7:0] ? $signed(regsB_82_re) : $signed(_GEN_8281); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8283 = 8'h31 == _T_31[7:0] ? $signed(regsB_92_re) : $signed(_GEN_8282); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8284 = 8'h32 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8283); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8285 = 8'h33 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8284); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8286 = 8'h34 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8285); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8287 = 8'h35 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8286); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8288 = 8'h36 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8287); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8289 = 8'h37 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8288); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8290 = 8'h38 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8289); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8291 = 8'h39 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8290); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8292 = 8'h3a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8291); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8293 = 8'h3b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8292); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8294 = 8'h3c == _T_31[7:0] ? $signed(regsB_3_re) : $signed(_GEN_8293); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8295 = 8'h3d == _T_31[7:0] ? $signed(regsB_13_re) : $signed(_GEN_8294); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8296 = 8'h3e == _T_31[7:0] ? $signed(regsB_23_re) : $signed(_GEN_8295); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8297 = 8'h3f == _T_31[7:0] ? $signed(regsB_33_re) : $signed(_GEN_8296); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8298 = 8'h40 == _T_31[7:0] ? $signed(regsB_43_re) : $signed(_GEN_8297); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8299 = 8'h41 == _T_31[7:0] ? $signed(regsB_53_re) : $signed(_GEN_8298); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8300 = 8'h42 == _T_31[7:0] ? $signed(regsB_63_re) : $signed(_GEN_8299); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8301 = 8'h43 == _T_31[7:0] ? $signed(regsB_73_re) : $signed(_GEN_8300); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8302 = 8'h44 == _T_31[7:0] ? $signed(regsB_83_re) : $signed(_GEN_8301); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8303 = 8'h45 == _T_31[7:0] ? $signed(regsB_93_re) : $signed(_GEN_8302); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8304 = 8'h46 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8303); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8305 = 8'h47 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8304); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8306 = 8'h48 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8305); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8307 = 8'h49 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8306); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8308 = 8'h4a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8307); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8309 = 8'h4b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8308); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8310 = 8'h4c == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8309); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8311 = 8'h4d == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8310); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8312 = 8'h4e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8311); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8313 = 8'h4f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8312); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8314 = 8'h50 == _T_31[7:0] ? $signed(regsB_4_re) : $signed(_GEN_8313); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8315 = 8'h51 == _T_31[7:0] ? $signed(regsB_14_re) : $signed(_GEN_8314); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8316 = 8'h52 == _T_31[7:0] ? $signed(regsB_24_re) : $signed(_GEN_8315); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8317 = 8'h53 == _T_31[7:0] ? $signed(regsB_34_re) : $signed(_GEN_8316); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8318 = 8'h54 == _T_31[7:0] ? $signed(regsB_44_re) : $signed(_GEN_8317); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8319 = 8'h55 == _T_31[7:0] ? $signed(regsB_54_re) : $signed(_GEN_8318); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8320 = 8'h56 == _T_31[7:0] ? $signed(regsB_64_re) : $signed(_GEN_8319); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8321 = 8'h57 == _T_31[7:0] ? $signed(regsB_74_re) : $signed(_GEN_8320); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8322 = 8'h58 == _T_31[7:0] ? $signed(regsB_84_re) : $signed(_GEN_8321); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8323 = 8'h59 == _T_31[7:0] ? $signed(regsB_94_re) : $signed(_GEN_8322); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8324 = 8'h5a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8323); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8325 = 8'h5b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8324); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8326 = 8'h5c == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8325); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8327 = 8'h5d == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8326); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8328 = 8'h5e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8327); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8329 = 8'h5f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8328); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8330 = 8'h60 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8329); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8331 = 8'h61 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8330); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8332 = 8'h62 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8331); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8333 = 8'h63 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8332); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8334 = 8'h64 == _T_31[7:0] ? $signed(regsB_5_re) : $signed(_GEN_8333); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8335 = 8'h65 == _T_31[7:0] ? $signed(regsB_15_re) : $signed(_GEN_8334); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8336 = 8'h66 == _T_31[7:0] ? $signed(regsB_25_re) : $signed(_GEN_8335); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8337 = 8'h67 == _T_31[7:0] ? $signed(regsB_35_re) : $signed(_GEN_8336); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8338 = 8'h68 == _T_31[7:0] ? $signed(regsB_45_re) : $signed(_GEN_8337); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8339 = 8'h69 == _T_31[7:0] ? $signed(regsB_55_re) : $signed(_GEN_8338); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8340 = 8'h6a == _T_31[7:0] ? $signed(regsB_65_re) : $signed(_GEN_8339); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8341 = 8'h6b == _T_31[7:0] ? $signed(regsB_75_re) : $signed(_GEN_8340); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8342 = 8'h6c == _T_31[7:0] ? $signed(regsB_85_re) : $signed(_GEN_8341); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8343 = 8'h6d == _T_31[7:0] ? $signed(regsB_95_re) : $signed(_GEN_8342); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8344 = 8'h6e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8343); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8345 = 8'h6f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8344); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8346 = 8'h70 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8345); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8347 = 8'h71 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8346); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8348 = 8'h72 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8347); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8349 = 8'h73 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8348); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8350 = 8'h74 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8349); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8351 = 8'h75 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8350); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8352 = 8'h76 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8351); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8353 = 8'h77 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8352); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8354 = 8'h78 == _T_31[7:0] ? $signed(regsB_6_re) : $signed(_GEN_8353); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8355 = 8'h79 == _T_31[7:0] ? $signed(regsB_16_re) : $signed(_GEN_8354); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8356 = 8'h7a == _T_31[7:0] ? $signed(regsB_26_re) : $signed(_GEN_8355); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8357 = 8'h7b == _T_31[7:0] ? $signed(regsB_36_re) : $signed(_GEN_8356); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8358 = 8'h7c == _T_31[7:0] ? $signed(regsB_46_re) : $signed(_GEN_8357); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8359 = 8'h7d == _T_31[7:0] ? $signed(regsB_56_re) : $signed(_GEN_8358); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8360 = 8'h7e == _T_31[7:0] ? $signed(regsB_66_re) : $signed(_GEN_8359); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8361 = 8'h7f == _T_31[7:0] ? $signed(regsB_76_re) : $signed(_GEN_8360); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8362 = 8'h80 == _T_31[7:0] ? $signed(regsB_86_re) : $signed(_GEN_8361); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8363 = 8'h81 == _T_31[7:0] ? $signed(regsB_96_re) : $signed(_GEN_8362); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8364 = 8'h82 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8363); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8365 = 8'h83 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8364); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8366 = 8'h84 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8365); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8367 = 8'h85 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8366); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8368 = 8'h86 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8367); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8369 = 8'h87 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8368); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8370 = 8'h88 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8369); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8371 = 8'h89 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8370); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8372 = 8'h8a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8371); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8373 = 8'h8b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8372); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8374 = 8'h8c == _T_31[7:0] ? $signed(regsB_7_re) : $signed(_GEN_8373); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8375 = 8'h8d == _T_31[7:0] ? $signed(regsB_17_re) : $signed(_GEN_8374); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8376 = 8'h8e == _T_31[7:0] ? $signed(regsB_27_re) : $signed(_GEN_8375); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8377 = 8'h8f == _T_31[7:0] ? $signed(regsB_37_re) : $signed(_GEN_8376); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8378 = 8'h90 == _T_31[7:0] ? $signed(regsB_47_re) : $signed(_GEN_8377); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8379 = 8'h91 == _T_31[7:0] ? $signed(regsB_57_re) : $signed(_GEN_8378); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8380 = 8'h92 == _T_31[7:0] ? $signed(regsB_67_re) : $signed(_GEN_8379); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8381 = 8'h93 == _T_31[7:0] ? $signed(regsB_77_re) : $signed(_GEN_8380); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8382 = 8'h94 == _T_31[7:0] ? $signed(regsB_87_re) : $signed(_GEN_8381); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8383 = 8'h95 == _T_31[7:0] ? $signed(regsB_97_re) : $signed(_GEN_8382); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8384 = 8'h96 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8383); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8385 = 8'h97 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8384); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8386 = 8'h98 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8385); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8387 = 8'h99 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8386); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8388 = 8'h9a == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8387); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8389 = 8'h9b == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8388); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8390 = 8'h9c == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8389); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8391 = 8'h9d == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8390); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8392 = 8'h9e == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8391); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8393 = 8'h9f == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8392); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8394 = 8'ha0 == _T_31[7:0] ? $signed(regsB_8_re) : $signed(_GEN_8393); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8395 = 8'ha1 == _T_31[7:0] ? $signed(regsB_18_re) : $signed(_GEN_8394); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8396 = 8'ha2 == _T_31[7:0] ? $signed(regsB_28_re) : $signed(_GEN_8395); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8397 = 8'ha3 == _T_31[7:0] ? $signed(regsB_38_re) : $signed(_GEN_8396); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8398 = 8'ha4 == _T_31[7:0] ? $signed(regsB_48_re) : $signed(_GEN_8397); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8399 = 8'ha5 == _T_31[7:0] ? $signed(regsB_58_re) : $signed(_GEN_8398); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8400 = 8'ha6 == _T_31[7:0] ? $signed(regsB_68_re) : $signed(_GEN_8399); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8401 = 8'ha7 == _T_31[7:0] ? $signed(regsB_78_re) : $signed(_GEN_8400); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8402 = 8'ha8 == _T_31[7:0] ? $signed(regsB_88_re) : $signed(_GEN_8401); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8403 = 8'ha9 == _T_31[7:0] ? $signed(regsB_98_re) : $signed(_GEN_8402); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8404 = 8'haa == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8403); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8405 = 8'hab == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8404); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8406 = 8'hac == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8405); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8407 = 8'had == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8406); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8408 = 8'hae == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8407); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8409 = 8'haf == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8408); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8410 = 8'hb0 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8409); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8411 = 8'hb1 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8410); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8412 = 8'hb2 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8411); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8413 = 8'hb3 == _T_31[7:0] ? $signed(32'sh0) : $signed(_GEN_8412); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8414 = 8'hb4 == _T_31[7:0] ? $signed(regsB_9_re) : $signed(_GEN_8413); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8415 = 8'hb5 == _T_31[7:0] ? $signed(regsB_19_re) : $signed(_GEN_8414); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8416 = 8'hb6 == _T_31[7:0] ? $signed(regsB_29_re) : $signed(_GEN_8415); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8417 = 8'hb7 == _T_31[7:0] ? $signed(regsB_39_re) : $signed(_GEN_8416); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8418 = 8'hb8 == _T_31[7:0] ? $signed(regsB_49_re) : $signed(_GEN_8417); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8419 = 8'hb9 == _T_31[7:0] ? $signed(regsB_59_re) : $signed(_GEN_8418); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8420 = 8'hba == _T_31[7:0] ? $signed(regsB_69_re) : $signed(_GEN_8419); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8421 = 8'hbb == _T_31[7:0] ? $signed(regsB_79_re) : $signed(_GEN_8420); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8422 = 8'hbc == _T_31[7:0] ? $signed(regsB_89_re) : $signed(_GEN_8421); // @[Matrix_Mul_V1.scala 162:{19,19}]
  wire [31:0] _GEN_8423 = 8'hbd == _T_31[7:0] ? $signed(regsB_99_re) : $signed(_GEN_8422); // @[Matrix_Mul_V1.scala 162:{19,19}]
  PE PE ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_clock),
    .io_reset(PE_io_reset),
    .io_in_x_re(PE_io_in_x_re),
    .io_in_x_im(PE_io_in_x_im),
    .io_in_y_re(PE_io_in_y_re),
    .io_in_y_im(PE_io_in_y_im),
    .io_out_pe_re(PE_io_out_pe_re),
    .io_out_pe_im(PE_io_out_pe_im),
    .io_out_x_re(PE_io_out_x_re),
    .io_out_x_im(PE_io_out_x_im),
    .io_out_y_re(PE_io_out_y_re),
    .io_out_y_im(PE_io_out_y_im)
  );
  PE PE_1 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_1_clock),
    .io_reset(PE_1_io_reset),
    .io_in_x_re(PE_1_io_in_x_re),
    .io_in_x_im(PE_1_io_in_x_im),
    .io_in_y_re(PE_1_io_in_y_re),
    .io_in_y_im(PE_1_io_in_y_im),
    .io_out_pe_re(PE_1_io_out_pe_re),
    .io_out_pe_im(PE_1_io_out_pe_im),
    .io_out_x_re(PE_1_io_out_x_re),
    .io_out_x_im(PE_1_io_out_x_im),
    .io_out_y_re(PE_1_io_out_y_re),
    .io_out_y_im(PE_1_io_out_y_im)
  );
  PE PE_2 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_2_clock),
    .io_reset(PE_2_io_reset),
    .io_in_x_re(PE_2_io_in_x_re),
    .io_in_x_im(PE_2_io_in_x_im),
    .io_in_y_re(PE_2_io_in_y_re),
    .io_in_y_im(PE_2_io_in_y_im),
    .io_out_pe_re(PE_2_io_out_pe_re),
    .io_out_pe_im(PE_2_io_out_pe_im),
    .io_out_x_re(PE_2_io_out_x_re),
    .io_out_x_im(PE_2_io_out_x_im),
    .io_out_y_re(PE_2_io_out_y_re),
    .io_out_y_im(PE_2_io_out_y_im)
  );
  PE PE_3 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_3_clock),
    .io_reset(PE_3_io_reset),
    .io_in_x_re(PE_3_io_in_x_re),
    .io_in_x_im(PE_3_io_in_x_im),
    .io_in_y_re(PE_3_io_in_y_re),
    .io_in_y_im(PE_3_io_in_y_im),
    .io_out_pe_re(PE_3_io_out_pe_re),
    .io_out_pe_im(PE_3_io_out_pe_im),
    .io_out_x_re(PE_3_io_out_x_re),
    .io_out_x_im(PE_3_io_out_x_im),
    .io_out_y_re(PE_3_io_out_y_re),
    .io_out_y_im(PE_3_io_out_y_im)
  );
  PE PE_4 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_4_clock),
    .io_reset(PE_4_io_reset),
    .io_in_x_re(PE_4_io_in_x_re),
    .io_in_x_im(PE_4_io_in_x_im),
    .io_in_y_re(PE_4_io_in_y_re),
    .io_in_y_im(PE_4_io_in_y_im),
    .io_out_pe_re(PE_4_io_out_pe_re),
    .io_out_pe_im(PE_4_io_out_pe_im),
    .io_out_x_re(PE_4_io_out_x_re),
    .io_out_x_im(PE_4_io_out_x_im),
    .io_out_y_re(PE_4_io_out_y_re),
    .io_out_y_im(PE_4_io_out_y_im)
  );
  PE PE_5 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_5_clock),
    .io_reset(PE_5_io_reset),
    .io_in_x_re(PE_5_io_in_x_re),
    .io_in_x_im(PE_5_io_in_x_im),
    .io_in_y_re(PE_5_io_in_y_re),
    .io_in_y_im(PE_5_io_in_y_im),
    .io_out_pe_re(PE_5_io_out_pe_re),
    .io_out_pe_im(PE_5_io_out_pe_im),
    .io_out_x_re(PE_5_io_out_x_re),
    .io_out_x_im(PE_5_io_out_x_im),
    .io_out_y_re(PE_5_io_out_y_re),
    .io_out_y_im(PE_5_io_out_y_im)
  );
  PE PE_6 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_6_clock),
    .io_reset(PE_6_io_reset),
    .io_in_x_re(PE_6_io_in_x_re),
    .io_in_x_im(PE_6_io_in_x_im),
    .io_in_y_re(PE_6_io_in_y_re),
    .io_in_y_im(PE_6_io_in_y_im),
    .io_out_pe_re(PE_6_io_out_pe_re),
    .io_out_pe_im(PE_6_io_out_pe_im),
    .io_out_x_re(PE_6_io_out_x_re),
    .io_out_x_im(PE_6_io_out_x_im),
    .io_out_y_re(PE_6_io_out_y_re),
    .io_out_y_im(PE_6_io_out_y_im)
  );
  PE PE_7 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_7_clock),
    .io_reset(PE_7_io_reset),
    .io_in_x_re(PE_7_io_in_x_re),
    .io_in_x_im(PE_7_io_in_x_im),
    .io_in_y_re(PE_7_io_in_y_re),
    .io_in_y_im(PE_7_io_in_y_im),
    .io_out_pe_re(PE_7_io_out_pe_re),
    .io_out_pe_im(PE_7_io_out_pe_im),
    .io_out_x_re(PE_7_io_out_x_re),
    .io_out_x_im(PE_7_io_out_x_im),
    .io_out_y_re(PE_7_io_out_y_re),
    .io_out_y_im(PE_7_io_out_y_im)
  );
  PE PE_8 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_8_clock),
    .io_reset(PE_8_io_reset),
    .io_in_x_re(PE_8_io_in_x_re),
    .io_in_x_im(PE_8_io_in_x_im),
    .io_in_y_re(PE_8_io_in_y_re),
    .io_in_y_im(PE_8_io_in_y_im),
    .io_out_pe_re(PE_8_io_out_pe_re),
    .io_out_pe_im(PE_8_io_out_pe_im),
    .io_out_x_re(PE_8_io_out_x_re),
    .io_out_x_im(PE_8_io_out_x_im),
    .io_out_y_re(PE_8_io_out_y_re),
    .io_out_y_im(PE_8_io_out_y_im)
  );
  PE PE_9 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_9_clock),
    .io_reset(PE_9_io_reset),
    .io_in_x_re(PE_9_io_in_x_re),
    .io_in_x_im(PE_9_io_in_x_im),
    .io_in_y_re(PE_9_io_in_y_re),
    .io_in_y_im(PE_9_io_in_y_im),
    .io_out_pe_re(PE_9_io_out_pe_re),
    .io_out_pe_im(PE_9_io_out_pe_im),
    .io_out_x_re(PE_9_io_out_x_re),
    .io_out_x_im(PE_9_io_out_x_im),
    .io_out_y_re(PE_9_io_out_y_re),
    .io_out_y_im(PE_9_io_out_y_im)
  );
  PE PE_10 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_10_clock),
    .io_reset(PE_10_io_reset),
    .io_in_x_re(PE_10_io_in_x_re),
    .io_in_x_im(PE_10_io_in_x_im),
    .io_in_y_re(PE_10_io_in_y_re),
    .io_in_y_im(PE_10_io_in_y_im),
    .io_out_pe_re(PE_10_io_out_pe_re),
    .io_out_pe_im(PE_10_io_out_pe_im),
    .io_out_x_re(PE_10_io_out_x_re),
    .io_out_x_im(PE_10_io_out_x_im),
    .io_out_y_re(PE_10_io_out_y_re),
    .io_out_y_im(PE_10_io_out_y_im)
  );
  PE PE_11 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_11_clock),
    .io_reset(PE_11_io_reset),
    .io_in_x_re(PE_11_io_in_x_re),
    .io_in_x_im(PE_11_io_in_x_im),
    .io_in_y_re(PE_11_io_in_y_re),
    .io_in_y_im(PE_11_io_in_y_im),
    .io_out_pe_re(PE_11_io_out_pe_re),
    .io_out_pe_im(PE_11_io_out_pe_im),
    .io_out_x_re(PE_11_io_out_x_re),
    .io_out_x_im(PE_11_io_out_x_im),
    .io_out_y_re(PE_11_io_out_y_re),
    .io_out_y_im(PE_11_io_out_y_im)
  );
  PE PE_12 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_12_clock),
    .io_reset(PE_12_io_reset),
    .io_in_x_re(PE_12_io_in_x_re),
    .io_in_x_im(PE_12_io_in_x_im),
    .io_in_y_re(PE_12_io_in_y_re),
    .io_in_y_im(PE_12_io_in_y_im),
    .io_out_pe_re(PE_12_io_out_pe_re),
    .io_out_pe_im(PE_12_io_out_pe_im),
    .io_out_x_re(PE_12_io_out_x_re),
    .io_out_x_im(PE_12_io_out_x_im),
    .io_out_y_re(PE_12_io_out_y_re),
    .io_out_y_im(PE_12_io_out_y_im)
  );
  PE PE_13 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_13_clock),
    .io_reset(PE_13_io_reset),
    .io_in_x_re(PE_13_io_in_x_re),
    .io_in_x_im(PE_13_io_in_x_im),
    .io_in_y_re(PE_13_io_in_y_re),
    .io_in_y_im(PE_13_io_in_y_im),
    .io_out_pe_re(PE_13_io_out_pe_re),
    .io_out_pe_im(PE_13_io_out_pe_im),
    .io_out_x_re(PE_13_io_out_x_re),
    .io_out_x_im(PE_13_io_out_x_im),
    .io_out_y_re(PE_13_io_out_y_re),
    .io_out_y_im(PE_13_io_out_y_im)
  );
  PE PE_14 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_14_clock),
    .io_reset(PE_14_io_reset),
    .io_in_x_re(PE_14_io_in_x_re),
    .io_in_x_im(PE_14_io_in_x_im),
    .io_in_y_re(PE_14_io_in_y_re),
    .io_in_y_im(PE_14_io_in_y_im),
    .io_out_pe_re(PE_14_io_out_pe_re),
    .io_out_pe_im(PE_14_io_out_pe_im),
    .io_out_x_re(PE_14_io_out_x_re),
    .io_out_x_im(PE_14_io_out_x_im),
    .io_out_y_re(PE_14_io_out_y_re),
    .io_out_y_im(PE_14_io_out_y_im)
  );
  PE PE_15 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_15_clock),
    .io_reset(PE_15_io_reset),
    .io_in_x_re(PE_15_io_in_x_re),
    .io_in_x_im(PE_15_io_in_x_im),
    .io_in_y_re(PE_15_io_in_y_re),
    .io_in_y_im(PE_15_io_in_y_im),
    .io_out_pe_re(PE_15_io_out_pe_re),
    .io_out_pe_im(PE_15_io_out_pe_im),
    .io_out_x_re(PE_15_io_out_x_re),
    .io_out_x_im(PE_15_io_out_x_im),
    .io_out_y_re(PE_15_io_out_y_re),
    .io_out_y_im(PE_15_io_out_y_im)
  );
  PE PE_16 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_16_clock),
    .io_reset(PE_16_io_reset),
    .io_in_x_re(PE_16_io_in_x_re),
    .io_in_x_im(PE_16_io_in_x_im),
    .io_in_y_re(PE_16_io_in_y_re),
    .io_in_y_im(PE_16_io_in_y_im),
    .io_out_pe_re(PE_16_io_out_pe_re),
    .io_out_pe_im(PE_16_io_out_pe_im),
    .io_out_x_re(PE_16_io_out_x_re),
    .io_out_x_im(PE_16_io_out_x_im),
    .io_out_y_re(PE_16_io_out_y_re),
    .io_out_y_im(PE_16_io_out_y_im)
  );
  PE PE_17 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_17_clock),
    .io_reset(PE_17_io_reset),
    .io_in_x_re(PE_17_io_in_x_re),
    .io_in_x_im(PE_17_io_in_x_im),
    .io_in_y_re(PE_17_io_in_y_re),
    .io_in_y_im(PE_17_io_in_y_im),
    .io_out_pe_re(PE_17_io_out_pe_re),
    .io_out_pe_im(PE_17_io_out_pe_im),
    .io_out_x_re(PE_17_io_out_x_re),
    .io_out_x_im(PE_17_io_out_x_im),
    .io_out_y_re(PE_17_io_out_y_re),
    .io_out_y_im(PE_17_io_out_y_im)
  );
  PE PE_18 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_18_clock),
    .io_reset(PE_18_io_reset),
    .io_in_x_re(PE_18_io_in_x_re),
    .io_in_x_im(PE_18_io_in_x_im),
    .io_in_y_re(PE_18_io_in_y_re),
    .io_in_y_im(PE_18_io_in_y_im),
    .io_out_pe_re(PE_18_io_out_pe_re),
    .io_out_pe_im(PE_18_io_out_pe_im),
    .io_out_x_re(PE_18_io_out_x_re),
    .io_out_x_im(PE_18_io_out_x_im),
    .io_out_y_re(PE_18_io_out_y_re),
    .io_out_y_im(PE_18_io_out_y_im)
  );
  PE PE_19 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_19_clock),
    .io_reset(PE_19_io_reset),
    .io_in_x_re(PE_19_io_in_x_re),
    .io_in_x_im(PE_19_io_in_x_im),
    .io_in_y_re(PE_19_io_in_y_re),
    .io_in_y_im(PE_19_io_in_y_im),
    .io_out_pe_re(PE_19_io_out_pe_re),
    .io_out_pe_im(PE_19_io_out_pe_im),
    .io_out_x_re(PE_19_io_out_x_re),
    .io_out_x_im(PE_19_io_out_x_im),
    .io_out_y_re(PE_19_io_out_y_re),
    .io_out_y_im(PE_19_io_out_y_im)
  );
  PE PE_20 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_20_clock),
    .io_reset(PE_20_io_reset),
    .io_in_x_re(PE_20_io_in_x_re),
    .io_in_x_im(PE_20_io_in_x_im),
    .io_in_y_re(PE_20_io_in_y_re),
    .io_in_y_im(PE_20_io_in_y_im),
    .io_out_pe_re(PE_20_io_out_pe_re),
    .io_out_pe_im(PE_20_io_out_pe_im),
    .io_out_x_re(PE_20_io_out_x_re),
    .io_out_x_im(PE_20_io_out_x_im),
    .io_out_y_re(PE_20_io_out_y_re),
    .io_out_y_im(PE_20_io_out_y_im)
  );
  PE PE_21 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_21_clock),
    .io_reset(PE_21_io_reset),
    .io_in_x_re(PE_21_io_in_x_re),
    .io_in_x_im(PE_21_io_in_x_im),
    .io_in_y_re(PE_21_io_in_y_re),
    .io_in_y_im(PE_21_io_in_y_im),
    .io_out_pe_re(PE_21_io_out_pe_re),
    .io_out_pe_im(PE_21_io_out_pe_im),
    .io_out_x_re(PE_21_io_out_x_re),
    .io_out_x_im(PE_21_io_out_x_im),
    .io_out_y_re(PE_21_io_out_y_re),
    .io_out_y_im(PE_21_io_out_y_im)
  );
  PE PE_22 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_22_clock),
    .io_reset(PE_22_io_reset),
    .io_in_x_re(PE_22_io_in_x_re),
    .io_in_x_im(PE_22_io_in_x_im),
    .io_in_y_re(PE_22_io_in_y_re),
    .io_in_y_im(PE_22_io_in_y_im),
    .io_out_pe_re(PE_22_io_out_pe_re),
    .io_out_pe_im(PE_22_io_out_pe_im),
    .io_out_x_re(PE_22_io_out_x_re),
    .io_out_x_im(PE_22_io_out_x_im),
    .io_out_y_re(PE_22_io_out_y_re),
    .io_out_y_im(PE_22_io_out_y_im)
  );
  PE PE_23 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_23_clock),
    .io_reset(PE_23_io_reset),
    .io_in_x_re(PE_23_io_in_x_re),
    .io_in_x_im(PE_23_io_in_x_im),
    .io_in_y_re(PE_23_io_in_y_re),
    .io_in_y_im(PE_23_io_in_y_im),
    .io_out_pe_re(PE_23_io_out_pe_re),
    .io_out_pe_im(PE_23_io_out_pe_im),
    .io_out_x_re(PE_23_io_out_x_re),
    .io_out_x_im(PE_23_io_out_x_im),
    .io_out_y_re(PE_23_io_out_y_re),
    .io_out_y_im(PE_23_io_out_y_im)
  );
  PE PE_24 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_24_clock),
    .io_reset(PE_24_io_reset),
    .io_in_x_re(PE_24_io_in_x_re),
    .io_in_x_im(PE_24_io_in_x_im),
    .io_in_y_re(PE_24_io_in_y_re),
    .io_in_y_im(PE_24_io_in_y_im),
    .io_out_pe_re(PE_24_io_out_pe_re),
    .io_out_pe_im(PE_24_io_out_pe_im),
    .io_out_x_re(PE_24_io_out_x_re),
    .io_out_x_im(PE_24_io_out_x_im),
    .io_out_y_re(PE_24_io_out_y_re),
    .io_out_y_im(PE_24_io_out_y_im)
  );
  PE PE_25 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_25_clock),
    .io_reset(PE_25_io_reset),
    .io_in_x_re(PE_25_io_in_x_re),
    .io_in_x_im(PE_25_io_in_x_im),
    .io_in_y_re(PE_25_io_in_y_re),
    .io_in_y_im(PE_25_io_in_y_im),
    .io_out_pe_re(PE_25_io_out_pe_re),
    .io_out_pe_im(PE_25_io_out_pe_im),
    .io_out_x_re(PE_25_io_out_x_re),
    .io_out_x_im(PE_25_io_out_x_im),
    .io_out_y_re(PE_25_io_out_y_re),
    .io_out_y_im(PE_25_io_out_y_im)
  );
  PE PE_26 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_26_clock),
    .io_reset(PE_26_io_reset),
    .io_in_x_re(PE_26_io_in_x_re),
    .io_in_x_im(PE_26_io_in_x_im),
    .io_in_y_re(PE_26_io_in_y_re),
    .io_in_y_im(PE_26_io_in_y_im),
    .io_out_pe_re(PE_26_io_out_pe_re),
    .io_out_pe_im(PE_26_io_out_pe_im),
    .io_out_x_re(PE_26_io_out_x_re),
    .io_out_x_im(PE_26_io_out_x_im),
    .io_out_y_re(PE_26_io_out_y_re),
    .io_out_y_im(PE_26_io_out_y_im)
  );
  PE PE_27 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_27_clock),
    .io_reset(PE_27_io_reset),
    .io_in_x_re(PE_27_io_in_x_re),
    .io_in_x_im(PE_27_io_in_x_im),
    .io_in_y_re(PE_27_io_in_y_re),
    .io_in_y_im(PE_27_io_in_y_im),
    .io_out_pe_re(PE_27_io_out_pe_re),
    .io_out_pe_im(PE_27_io_out_pe_im),
    .io_out_x_re(PE_27_io_out_x_re),
    .io_out_x_im(PE_27_io_out_x_im),
    .io_out_y_re(PE_27_io_out_y_re),
    .io_out_y_im(PE_27_io_out_y_im)
  );
  PE PE_28 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_28_clock),
    .io_reset(PE_28_io_reset),
    .io_in_x_re(PE_28_io_in_x_re),
    .io_in_x_im(PE_28_io_in_x_im),
    .io_in_y_re(PE_28_io_in_y_re),
    .io_in_y_im(PE_28_io_in_y_im),
    .io_out_pe_re(PE_28_io_out_pe_re),
    .io_out_pe_im(PE_28_io_out_pe_im),
    .io_out_x_re(PE_28_io_out_x_re),
    .io_out_x_im(PE_28_io_out_x_im),
    .io_out_y_re(PE_28_io_out_y_re),
    .io_out_y_im(PE_28_io_out_y_im)
  );
  PE PE_29 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_29_clock),
    .io_reset(PE_29_io_reset),
    .io_in_x_re(PE_29_io_in_x_re),
    .io_in_x_im(PE_29_io_in_x_im),
    .io_in_y_re(PE_29_io_in_y_re),
    .io_in_y_im(PE_29_io_in_y_im),
    .io_out_pe_re(PE_29_io_out_pe_re),
    .io_out_pe_im(PE_29_io_out_pe_im),
    .io_out_x_re(PE_29_io_out_x_re),
    .io_out_x_im(PE_29_io_out_x_im),
    .io_out_y_re(PE_29_io_out_y_re),
    .io_out_y_im(PE_29_io_out_y_im)
  );
  PE PE_30 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_30_clock),
    .io_reset(PE_30_io_reset),
    .io_in_x_re(PE_30_io_in_x_re),
    .io_in_x_im(PE_30_io_in_x_im),
    .io_in_y_re(PE_30_io_in_y_re),
    .io_in_y_im(PE_30_io_in_y_im),
    .io_out_pe_re(PE_30_io_out_pe_re),
    .io_out_pe_im(PE_30_io_out_pe_im),
    .io_out_x_re(PE_30_io_out_x_re),
    .io_out_x_im(PE_30_io_out_x_im),
    .io_out_y_re(PE_30_io_out_y_re),
    .io_out_y_im(PE_30_io_out_y_im)
  );
  PE PE_31 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_31_clock),
    .io_reset(PE_31_io_reset),
    .io_in_x_re(PE_31_io_in_x_re),
    .io_in_x_im(PE_31_io_in_x_im),
    .io_in_y_re(PE_31_io_in_y_re),
    .io_in_y_im(PE_31_io_in_y_im),
    .io_out_pe_re(PE_31_io_out_pe_re),
    .io_out_pe_im(PE_31_io_out_pe_im),
    .io_out_x_re(PE_31_io_out_x_re),
    .io_out_x_im(PE_31_io_out_x_im),
    .io_out_y_re(PE_31_io_out_y_re),
    .io_out_y_im(PE_31_io_out_y_im)
  );
  PE PE_32 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_32_clock),
    .io_reset(PE_32_io_reset),
    .io_in_x_re(PE_32_io_in_x_re),
    .io_in_x_im(PE_32_io_in_x_im),
    .io_in_y_re(PE_32_io_in_y_re),
    .io_in_y_im(PE_32_io_in_y_im),
    .io_out_pe_re(PE_32_io_out_pe_re),
    .io_out_pe_im(PE_32_io_out_pe_im),
    .io_out_x_re(PE_32_io_out_x_re),
    .io_out_x_im(PE_32_io_out_x_im),
    .io_out_y_re(PE_32_io_out_y_re),
    .io_out_y_im(PE_32_io_out_y_im)
  );
  PE PE_33 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_33_clock),
    .io_reset(PE_33_io_reset),
    .io_in_x_re(PE_33_io_in_x_re),
    .io_in_x_im(PE_33_io_in_x_im),
    .io_in_y_re(PE_33_io_in_y_re),
    .io_in_y_im(PE_33_io_in_y_im),
    .io_out_pe_re(PE_33_io_out_pe_re),
    .io_out_pe_im(PE_33_io_out_pe_im),
    .io_out_x_re(PE_33_io_out_x_re),
    .io_out_x_im(PE_33_io_out_x_im),
    .io_out_y_re(PE_33_io_out_y_re),
    .io_out_y_im(PE_33_io_out_y_im)
  );
  PE PE_34 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_34_clock),
    .io_reset(PE_34_io_reset),
    .io_in_x_re(PE_34_io_in_x_re),
    .io_in_x_im(PE_34_io_in_x_im),
    .io_in_y_re(PE_34_io_in_y_re),
    .io_in_y_im(PE_34_io_in_y_im),
    .io_out_pe_re(PE_34_io_out_pe_re),
    .io_out_pe_im(PE_34_io_out_pe_im),
    .io_out_x_re(PE_34_io_out_x_re),
    .io_out_x_im(PE_34_io_out_x_im),
    .io_out_y_re(PE_34_io_out_y_re),
    .io_out_y_im(PE_34_io_out_y_im)
  );
  PE PE_35 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_35_clock),
    .io_reset(PE_35_io_reset),
    .io_in_x_re(PE_35_io_in_x_re),
    .io_in_x_im(PE_35_io_in_x_im),
    .io_in_y_re(PE_35_io_in_y_re),
    .io_in_y_im(PE_35_io_in_y_im),
    .io_out_pe_re(PE_35_io_out_pe_re),
    .io_out_pe_im(PE_35_io_out_pe_im),
    .io_out_x_re(PE_35_io_out_x_re),
    .io_out_x_im(PE_35_io_out_x_im),
    .io_out_y_re(PE_35_io_out_y_re),
    .io_out_y_im(PE_35_io_out_y_im)
  );
  PE PE_36 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_36_clock),
    .io_reset(PE_36_io_reset),
    .io_in_x_re(PE_36_io_in_x_re),
    .io_in_x_im(PE_36_io_in_x_im),
    .io_in_y_re(PE_36_io_in_y_re),
    .io_in_y_im(PE_36_io_in_y_im),
    .io_out_pe_re(PE_36_io_out_pe_re),
    .io_out_pe_im(PE_36_io_out_pe_im),
    .io_out_x_re(PE_36_io_out_x_re),
    .io_out_x_im(PE_36_io_out_x_im),
    .io_out_y_re(PE_36_io_out_y_re),
    .io_out_y_im(PE_36_io_out_y_im)
  );
  PE PE_37 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_37_clock),
    .io_reset(PE_37_io_reset),
    .io_in_x_re(PE_37_io_in_x_re),
    .io_in_x_im(PE_37_io_in_x_im),
    .io_in_y_re(PE_37_io_in_y_re),
    .io_in_y_im(PE_37_io_in_y_im),
    .io_out_pe_re(PE_37_io_out_pe_re),
    .io_out_pe_im(PE_37_io_out_pe_im),
    .io_out_x_re(PE_37_io_out_x_re),
    .io_out_x_im(PE_37_io_out_x_im),
    .io_out_y_re(PE_37_io_out_y_re),
    .io_out_y_im(PE_37_io_out_y_im)
  );
  PE PE_38 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_38_clock),
    .io_reset(PE_38_io_reset),
    .io_in_x_re(PE_38_io_in_x_re),
    .io_in_x_im(PE_38_io_in_x_im),
    .io_in_y_re(PE_38_io_in_y_re),
    .io_in_y_im(PE_38_io_in_y_im),
    .io_out_pe_re(PE_38_io_out_pe_re),
    .io_out_pe_im(PE_38_io_out_pe_im),
    .io_out_x_re(PE_38_io_out_x_re),
    .io_out_x_im(PE_38_io_out_x_im),
    .io_out_y_re(PE_38_io_out_y_re),
    .io_out_y_im(PE_38_io_out_y_im)
  );
  PE PE_39 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_39_clock),
    .io_reset(PE_39_io_reset),
    .io_in_x_re(PE_39_io_in_x_re),
    .io_in_x_im(PE_39_io_in_x_im),
    .io_in_y_re(PE_39_io_in_y_re),
    .io_in_y_im(PE_39_io_in_y_im),
    .io_out_pe_re(PE_39_io_out_pe_re),
    .io_out_pe_im(PE_39_io_out_pe_im),
    .io_out_x_re(PE_39_io_out_x_re),
    .io_out_x_im(PE_39_io_out_x_im),
    .io_out_y_re(PE_39_io_out_y_re),
    .io_out_y_im(PE_39_io_out_y_im)
  );
  PE PE_40 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_40_clock),
    .io_reset(PE_40_io_reset),
    .io_in_x_re(PE_40_io_in_x_re),
    .io_in_x_im(PE_40_io_in_x_im),
    .io_in_y_re(PE_40_io_in_y_re),
    .io_in_y_im(PE_40_io_in_y_im),
    .io_out_pe_re(PE_40_io_out_pe_re),
    .io_out_pe_im(PE_40_io_out_pe_im),
    .io_out_x_re(PE_40_io_out_x_re),
    .io_out_x_im(PE_40_io_out_x_im),
    .io_out_y_re(PE_40_io_out_y_re),
    .io_out_y_im(PE_40_io_out_y_im)
  );
  PE PE_41 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_41_clock),
    .io_reset(PE_41_io_reset),
    .io_in_x_re(PE_41_io_in_x_re),
    .io_in_x_im(PE_41_io_in_x_im),
    .io_in_y_re(PE_41_io_in_y_re),
    .io_in_y_im(PE_41_io_in_y_im),
    .io_out_pe_re(PE_41_io_out_pe_re),
    .io_out_pe_im(PE_41_io_out_pe_im),
    .io_out_x_re(PE_41_io_out_x_re),
    .io_out_x_im(PE_41_io_out_x_im),
    .io_out_y_re(PE_41_io_out_y_re),
    .io_out_y_im(PE_41_io_out_y_im)
  );
  PE PE_42 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_42_clock),
    .io_reset(PE_42_io_reset),
    .io_in_x_re(PE_42_io_in_x_re),
    .io_in_x_im(PE_42_io_in_x_im),
    .io_in_y_re(PE_42_io_in_y_re),
    .io_in_y_im(PE_42_io_in_y_im),
    .io_out_pe_re(PE_42_io_out_pe_re),
    .io_out_pe_im(PE_42_io_out_pe_im),
    .io_out_x_re(PE_42_io_out_x_re),
    .io_out_x_im(PE_42_io_out_x_im),
    .io_out_y_re(PE_42_io_out_y_re),
    .io_out_y_im(PE_42_io_out_y_im)
  );
  PE PE_43 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_43_clock),
    .io_reset(PE_43_io_reset),
    .io_in_x_re(PE_43_io_in_x_re),
    .io_in_x_im(PE_43_io_in_x_im),
    .io_in_y_re(PE_43_io_in_y_re),
    .io_in_y_im(PE_43_io_in_y_im),
    .io_out_pe_re(PE_43_io_out_pe_re),
    .io_out_pe_im(PE_43_io_out_pe_im),
    .io_out_x_re(PE_43_io_out_x_re),
    .io_out_x_im(PE_43_io_out_x_im),
    .io_out_y_re(PE_43_io_out_y_re),
    .io_out_y_im(PE_43_io_out_y_im)
  );
  PE PE_44 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_44_clock),
    .io_reset(PE_44_io_reset),
    .io_in_x_re(PE_44_io_in_x_re),
    .io_in_x_im(PE_44_io_in_x_im),
    .io_in_y_re(PE_44_io_in_y_re),
    .io_in_y_im(PE_44_io_in_y_im),
    .io_out_pe_re(PE_44_io_out_pe_re),
    .io_out_pe_im(PE_44_io_out_pe_im),
    .io_out_x_re(PE_44_io_out_x_re),
    .io_out_x_im(PE_44_io_out_x_im),
    .io_out_y_re(PE_44_io_out_y_re),
    .io_out_y_im(PE_44_io_out_y_im)
  );
  PE PE_45 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_45_clock),
    .io_reset(PE_45_io_reset),
    .io_in_x_re(PE_45_io_in_x_re),
    .io_in_x_im(PE_45_io_in_x_im),
    .io_in_y_re(PE_45_io_in_y_re),
    .io_in_y_im(PE_45_io_in_y_im),
    .io_out_pe_re(PE_45_io_out_pe_re),
    .io_out_pe_im(PE_45_io_out_pe_im),
    .io_out_x_re(PE_45_io_out_x_re),
    .io_out_x_im(PE_45_io_out_x_im),
    .io_out_y_re(PE_45_io_out_y_re),
    .io_out_y_im(PE_45_io_out_y_im)
  );
  PE PE_46 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_46_clock),
    .io_reset(PE_46_io_reset),
    .io_in_x_re(PE_46_io_in_x_re),
    .io_in_x_im(PE_46_io_in_x_im),
    .io_in_y_re(PE_46_io_in_y_re),
    .io_in_y_im(PE_46_io_in_y_im),
    .io_out_pe_re(PE_46_io_out_pe_re),
    .io_out_pe_im(PE_46_io_out_pe_im),
    .io_out_x_re(PE_46_io_out_x_re),
    .io_out_x_im(PE_46_io_out_x_im),
    .io_out_y_re(PE_46_io_out_y_re),
    .io_out_y_im(PE_46_io_out_y_im)
  );
  PE PE_47 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_47_clock),
    .io_reset(PE_47_io_reset),
    .io_in_x_re(PE_47_io_in_x_re),
    .io_in_x_im(PE_47_io_in_x_im),
    .io_in_y_re(PE_47_io_in_y_re),
    .io_in_y_im(PE_47_io_in_y_im),
    .io_out_pe_re(PE_47_io_out_pe_re),
    .io_out_pe_im(PE_47_io_out_pe_im),
    .io_out_x_re(PE_47_io_out_x_re),
    .io_out_x_im(PE_47_io_out_x_im),
    .io_out_y_re(PE_47_io_out_y_re),
    .io_out_y_im(PE_47_io_out_y_im)
  );
  PE PE_48 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_48_clock),
    .io_reset(PE_48_io_reset),
    .io_in_x_re(PE_48_io_in_x_re),
    .io_in_x_im(PE_48_io_in_x_im),
    .io_in_y_re(PE_48_io_in_y_re),
    .io_in_y_im(PE_48_io_in_y_im),
    .io_out_pe_re(PE_48_io_out_pe_re),
    .io_out_pe_im(PE_48_io_out_pe_im),
    .io_out_x_re(PE_48_io_out_x_re),
    .io_out_x_im(PE_48_io_out_x_im),
    .io_out_y_re(PE_48_io_out_y_re),
    .io_out_y_im(PE_48_io_out_y_im)
  );
  PE PE_49 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_49_clock),
    .io_reset(PE_49_io_reset),
    .io_in_x_re(PE_49_io_in_x_re),
    .io_in_x_im(PE_49_io_in_x_im),
    .io_in_y_re(PE_49_io_in_y_re),
    .io_in_y_im(PE_49_io_in_y_im),
    .io_out_pe_re(PE_49_io_out_pe_re),
    .io_out_pe_im(PE_49_io_out_pe_im),
    .io_out_x_re(PE_49_io_out_x_re),
    .io_out_x_im(PE_49_io_out_x_im),
    .io_out_y_re(PE_49_io_out_y_re),
    .io_out_y_im(PE_49_io_out_y_im)
  );
  PE PE_50 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_50_clock),
    .io_reset(PE_50_io_reset),
    .io_in_x_re(PE_50_io_in_x_re),
    .io_in_x_im(PE_50_io_in_x_im),
    .io_in_y_re(PE_50_io_in_y_re),
    .io_in_y_im(PE_50_io_in_y_im),
    .io_out_pe_re(PE_50_io_out_pe_re),
    .io_out_pe_im(PE_50_io_out_pe_im),
    .io_out_x_re(PE_50_io_out_x_re),
    .io_out_x_im(PE_50_io_out_x_im),
    .io_out_y_re(PE_50_io_out_y_re),
    .io_out_y_im(PE_50_io_out_y_im)
  );
  PE PE_51 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_51_clock),
    .io_reset(PE_51_io_reset),
    .io_in_x_re(PE_51_io_in_x_re),
    .io_in_x_im(PE_51_io_in_x_im),
    .io_in_y_re(PE_51_io_in_y_re),
    .io_in_y_im(PE_51_io_in_y_im),
    .io_out_pe_re(PE_51_io_out_pe_re),
    .io_out_pe_im(PE_51_io_out_pe_im),
    .io_out_x_re(PE_51_io_out_x_re),
    .io_out_x_im(PE_51_io_out_x_im),
    .io_out_y_re(PE_51_io_out_y_re),
    .io_out_y_im(PE_51_io_out_y_im)
  );
  PE PE_52 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_52_clock),
    .io_reset(PE_52_io_reset),
    .io_in_x_re(PE_52_io_in_x_re),
    .io_in_x_im(PE_52_io_in_x_im),
    .io_in_y_re(PE_52_io_in_y_re),
    .io_in_y_im(PE_52_io_in_y_im),
    .io_out_pe_re(PE_52_io_out_pe_re),
    .io_out_pe_im(PE_52_io_out_pe_im),
    .io_out_x_re(PE_52_io_out_x_re),
    .io_out_x_im(PE_52_io_out_x_im),
    .io_out_y_re(PE_52_io_out_y_re),
    .io_out_y_im(PE_52_io_out_y_im)
  );
  PE PE_53 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_53_clock),
    .io_reset(PE_53_io_reset),
    .io_in_x_re(PE_53_io_in_x_re),
    .io_in_x_im(PE_53_io_in_x_im),
    .io_in_y_re(PE_53_io_in_y_re),
    .io_in_y_im(PE_53_io_in_y_im),
    .io_out_pe_re(PE_53_io_out_pe_re),
    .io_out_pe_im(PE_53_io_out_pe_im),
    .io_out_x_re(PE_53_io_out_x_re),
    .io_out_x_im(PE_53_io_out_x_im),
    .io_out_y_re(PE_53_io_out_y_re),
    .io_out_y_im(PE_53_io_out_y_im)
  );
  PE PE_54 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_54_clock),
    .io_reset(PE_54_io_reset),
    .io_in_x_re(PE_54_io_in_x_re),
    .io_in_x_im(PE_54_io_in_x_im),
    .io_in_y_re(PE_54_io_in_y_re),
    .io_in_y_im(PE_54_io_in_y_im),
    .io_out_pe_re(PE_54_io_out_pe_re),
    .io_out_pe_im(PE_54_io_out_pe_im),
    .io_out_x_re(PE_54_io_out_x_re),
    .io_out_x_im(PE_54_io_out_x_im),
    .io_out_y_re(PE_54_io_out_y_re),
    .io_out_y_im(PE_54_io_out_y_im)
  );
  PE PE_55 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_55_clock),
    .io_reset(PE_55_io_reset),
    .io_in_x_re(PE_55_io_in_x_re),
    .io_in_x_im(PE_55_io_in_x_im),
    .io_in_y_re(PE_55_io_in_y_re),
    .io_in_y_im(PE_55_io_in_y_im),
    .io_out_pe_re(PE_55_io_out_pe_re),
    .io_out_pe_im(PE_55_io_out_pe_im),
    .io_out_x_re(PE_55_io_out_x_re),
    .io_out_x_im(PE_55_io_out_x_im),
    .io_out_y_re(PE_55_io_out_y_re),
    .io_out_y_im(PE_55_io_out_y_im)
  );
  PE PE_56 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_56_clock),
    .io_reset(PE_56_io_reset),
    .io_in_x_re(PE_56_io_in_x_re),
    .io_in_x_im(PE_56_io_in_x_im),
    .io_in_y_re(PE_56_io_in_y_re),
    .io_in_y_im(PE_56_io_in_y_im),
    .io_out_pe_re(PE_56_io_out_pe_re),
    .io_out_pe_im(PE_56_io_out_pe_im),
    .io_out_x_re(PE_56_io_out_x_re),
    .io_out_x_im(PE_56_io_out_x_im),
    .io_out_y_re(PE_56_io_out_y_re),
    .io_out_y_im(PE_56_io_out_y_im)
  );
  PE PE_57 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_57_clock),
    .io_reset(PE_57_io_reset),
    .io_in_x_re(PE_57_io_in_x_re),
    .io_in_x_im(PE_57_io_in_x_im),
    .io_in_y_re(PE_57_io_in_y_re),
    .io_in_y_im(PE_57_io_in_y_im),
    .io_out_pe_re(PE_57_io_out_pe_re),
    .io_out_pe_im(PE_57_io_out_pe_im),
    .io_out_x_re(PE_57_io_out_x_re),
    .io_out_x_im(PE_57_io_out_x_im),
    .io_out_y_re(PE_57_io_out_y_re),
    .io_out_y_im(PE_57_io_out_y_im)
  );
  PE PE_58 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_58_clock),
    .io_reset(PE_58_io_reset),
    .io_in_x_re(PE_58_io_in_x_re),
    .io_in_x_im(PE_58_io_in_x_im),
    .io_in_y_re(PE_58_io_in_y_re),
    .io_in_y_im(PE_58_io_in_y_im),
    .io_out_pe_re(PE_58_io_out_pe_re),
    .io_out_pe_im(PE_58_io_out_pe_im),
    .io_out_x_re(PE_58_io_out_x_re),
    .io_out_x_im(PE_58_io_out_x_im),
    .io_out_y_re(PE_58_io_out_y_re),
    .io_out_y_im(PE_58_io_out_y_im)
  );
  PE PE_59 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_59_clock),
    .io_reset(PE_59_io_reset),
    .io_in_x_re(PE_59_io_in_x_re),
    .io_in_x_im(PE_59_io_in_x_im),
    .io_in_y_re(PE_59_io_in_y_re),
    .io_in_y_im(PE_59_io_in_y_im),
    .io_out_pe_re(PE_59_io_out_pe_re),
    .io_out_pe_im(PE_59_io_out_pe_im),
    .io_out_x_re(PE_59_io_out_x_re),
    .io_out_x_im(PE_59_io_out_x_im),
    .io_out_y_re(PE_59_io_out_y_re),
    .io_out_y_im(PE_59_io_out_y_im)
  );
  PE PE_60 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_60_clock),
    .io_reset(PE_60_io_reset),
    .io_in_x_re(PE_60_io_in_x_re),
    .io_in_x_im(PE_60_io_in_x_im),
    .io_in_y_re(PE_60_io_in_y_re),
    .io_in_y_im(PE_60_io_in_y_im),
    .io_out_pe_re(PE_60_io_out_pe_re),
    .io_out_pe_im(PE_60_io_out_pe_im),
    .io_out_x_re(PE_60_io_out_x_re),
    .io_out_x_im(PE_60_io_out_x_im),
    .io_out_y_re(PE_60_io_out_y_re),
    .io_out_y_im(PE_60_io_out_y_im)
  );
  PE PE_61 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_61_clock),
    .io_reset(PE_61_io_reset),
    .io_in_x_re(PE_61_io_in_x_re),
    .io_in_x_im(PE_61_io_in_x_im),
    .io_in_y_re(PE_61_io_in_y_re),
    .io_in_y_im(PE_61_io_in_y_im),
    .io_out_pe_re(PE_61_io_out_pe_re),
    .io_out_pe_im(PE_61_io_out_pe_im),
    .io_out_x_re(PE_61_io_out_x_re),
    .io_out_x_im(PE_61_io_out_x_im),
    .io_out_y_re(PE_61_io_out_y_re),
    .io_out_y_im(PE_61_io_out_y_im)
  );
  PE PE_62 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_62_clock),
    .io_reset(PE_62_io_reset),
    .io_in_x_re(PE_62_io_in_x_re),
    .io_in_x_im(PE_62_io_in_x_im),
    .io_in_y_re(PE_62_io_in_y_re),
    .io_in_y_im(PE_62_io_in_y_im),
    .io_out_pe_re(PE_62_io_out_pe_re),
    .io_out_pe_im(PE_62_io_out_pe_im),
    .io_out_x_re(PE_62_io_out_x_re),
    .io_out_x_im(PE_62_io_out_x_im),
    .io_out_y_re(PE_62_io_out_y_re),
    .io_out_y_im(PE_62_io_out_y_im)
  );
  PE PE_63 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_63_clock),
    .io_reset(PE_63_io_reset),
    .io_in_x_re(PE_63_io_in_x_re),
    .io_in_x_im(PE_63_io_in_x_im),
    .io_in_y_re(PE_63_io_in_y_re),
    .io_in_y_im(PE_63_io_in_y_im),
    .io_out_pe_re(PE_63_io_out_pe_re),
    .io_out_pe_im(PE_63_io_out_pe_im),
    .io_out_x_re(PE_63_io_out_x_re),
    .io_out_x_im(PE_63_io_out_x_im),
    .io_out_y_re(PE_63_io_out_y_re),
    .io_out_y_im(PE_63_io_out_y_im)
  );
  PE PE_64 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_64_clock),
    .io_reset(PE_64_io_reset),
    .io_in_x_re(PE_64_io_in_x_re),
    .io_in_x_im(PE_64_io_in_x_im),
    .io_in_y_re(PE_64_io_in_y_re),
    .io_in_y_im(PE_64_io_in_y_im),
    .io_out_pe_re(PE_64_io_out_pe_re),
    .io_out_pe_im(PE_64_io_out_pe_im),
    .io_out_x_re(PE_64_io_out_x_re),
    .io_out_x_im(PE_64_io_out_x_im),
    .io_out_y_re(PE_64_io_out_y_re),
    .io_out_y_im(PE_64_io_out_y_im)
  );
  PE PE_65 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_65_clock),
    .io_reset(PE_65_io_reset),
    .io_in_x_re(PE_65_io_in_x_re),
    .io_in_x_im(PE_65_io_in_x_im),
    .io_in_y_re(PE_65_io_in_y_re),
    .io_in_y_im(PE_65_io_in_y_im),
    .io_out_pe_re(PE_65_io_out_pe_re),
    .io_out_pe_im(PE_65_io_out_pe_im),
    .io_out_x_re(PE_65_io_out_x_re),
    .io_out_x_im(PE_65_io_out_x_im),
    .io_out_y_re(PE_65_io_out_y_re),
    .io_out_y_im(PE_65_io_out_y_im)
  );
  PE PE_66 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_66_clock),
    .io_reset(PE_66_io_reset),
    .io_in_x_re(PE_66_io_in_x_re),
    .io_in_x_im(PE_66_io_in_x_im),
    .io_in_y_re(PE_66_io_in_y_re),
    .io_in_y_im(PE_66_io_in_y_im),
    .io_out_pe_re(PE_66_io_out_pe_re),
    .io_out_pe_im(PE_66_io_out_pe_im),
    .io_out_x_re(PE_66_io_out_x_re),
    .io_out_x_im(PE_66_io_out_x_im),
    .io_out_y_re(PE_66_io_out_y_re),
    .io_out_y_im(PE_66_io_out_y_im)
  );
  PE PE_67 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_67_clock),
    .io_reset(PE_67_io_reset),
    .io_in_x_re(PE_67_io_in_x_re),
    .io_in_x_im(PE_67_io_in_x_im),
    .io_in_y_re(PE_67_io_in_y_re),
    .io_in_y_im(PE_67_io_in_y_im),
    .io_out_pe_re(PE_67_io_out_pe_re),
    .io_out_pe_im(PE_67_io_out_pe_im),
    .io_out_x_re(PE_67_io_out_x_re),
    .io_out_x_im(PE_67_io_out_x_im),
    .io_out_y_re(PE_67_io_out_y_re),
    .io_out_y_im(PE_67_io_out_y_im)
  );
  PE PE_68 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_68_clock),
    .io_reset(PE_68_io_reset),
    .io_in_x_re(PE_68_io_in_x_re),
    .io_in_x_im(PE_68_io_in_x_im),
    .io_in_y_re(PE_68_io_in_y_re),
    .io_in_y_im(PE_68_io_in_y_im),
    .io_out_pe_re(PE_68_io_out_pe_re),
    .io_out_pe_im(PE_68_io_out_pe_im),
    .io_out_x_re(PE_68_io_out_x_re),
    .io_out_x_im(PE_68_io_out_x_im),
    .io_out_y_re(PE_68_io_out_y_re),
    .io_out_y_im(PE_68_io_out_y_im)
  );
  PE PE_69 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_69_clock),
    .io_reset(PE_69_io_reset),
    .io_in_x_re(PE_69_io_in_x_re),
    .io_in_x_im(PE_69_io_in_x_im),
    .io_in_y_re(PE_69_io_in_y_re),
    .io_in_y_im(PE_69_io_in_y_im),
    .io_out_pe_re(PE_69_io_out_pe_re),
    .io_out_pe_im(PE_69_io_out_pe_im),
    .io_out_x_re(PE_69_io_out_x_re),
    .io_out_x_im(PE_69_io_out_x_im),
    .io_out_y_re(PE_69_io_out_y_re),
    .io_out_y_im(PE_69_io_out_y_im)
  );
  PE PE_70 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_70_clock),
    .io_reset(PE_70_io_reset),
    .io_in_x_re(PE_70_io_in_x_re),
    .io_in_x_im(PE_70_io_in_x_im),
    .io_in_y_re(PE_70_io_in_y_re),
    .io_in_y_im(PE_70_io_in_y_im),
    .io_out_pe_re(PE_70_io_out_pe_re),
    .io_out_pe_im(PE_70_io_out_pe_im),
    .io_out_x_re(PE_70_io_out_x_re),
    .io_out_x_im(PE_70_io_out_x_im),
    .io_out_y_re(PE_70_io_out_y_re),
    .io_out_y_im(PE_70_io_out_y_im)
  );
  PE PE_71 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_71_clock),
    .io_reset(PE_71_io_reset),
    .io_in_x_re(PE_71_io_in_x_re),
    .io_in_x_im(PE_71_io_in_x_im),
    .io_in_y_re(PE_71_io_in_y_re),
    .io_in_y_im(PE_71_io_in_y_im),
    .io_out_pe_re(PE_71_io_out_pe_re),
    .io_out_pe_im(PE_71_io_out_pe_im),
    .io_out_x_re(PE_71_io_out_x_re),
    .io_out_x_im(PE_71_io_out_x_im),
    .io_out_y_re(PE_71_io_out_y_re),
    .io_out_y_im(PE_71_io_out_y_im)
  );
  PE PE_72 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_72_clock),
    .io_reset(PE_72_io_reset),
    .io_in_x_re(PE_72_io_in_x_re),
    .io_in_x_im(PE_72_io_in_x_im),
    .io_in_y_re(PE_72_io_in_y_re),
    .io_in_y_im(PE_72_io_in_y_im),
    .io_out_pe_re(PE_72_io_out_pe_re),
    .io_out_pe_im(PE_72_io_out_pe_im),
    .io_out_x_re(PE_72_io_out_x_re),
    .io_out_x_im(PE_72_io_out_x_im),
    .io_out_y_re(PE_72_io_out_y_re),
    .io_out_y_im(PE_72_io_out_y_im)
  );
  PE PE_73 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_73_clock),
    .io_reset(PE_73_io_reset),
    .io_in_x_re(PE_73_io_in_x_re),
    .io_in_x_im(PE_73_io_in_x_im),
    .io_in_y_re(PE_73_io_in_y_re),
    .io_in_y_im(PE_73_io_in_y_im),
    .io_out_pe_re(PE_73_io_out_pe_re),
    .io_out_pe_im(PE_73_io_out_pe_im),
    .io_out_x_re(PE_73_io_out_x_re),
    .io_out_x_im(PE_73_io_out_x_im),
    .io_out_y_re(PE_73_io_out_y_re),
    .io_out_y_im(PE_73_io_out_y_im)
  );
  PE PE_74 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_74_clock),
    .io_reset(PE_74_io_reset),
    .io_in_x_re(PE_74_io_in_x_re),
    .io_in_x_im(PE_74_io_in_x_im),
    .io_in_y_re(PE_74_io_in_y_re),
    .io_in_y_im(PE_74_io_in_y_im),
    .io_out_pe_re(PE_74_io_out_pe_re),
    .io_out_pe_im(PE_74_io_out_pe_im),
    .io_out_x_re(PE_74_io_out_x_re),
    .io_out_x_im(PE_74_io_out_x_im),
    .io_out_y_re(PE_74_io_out_y_re),
    .io_out_y_im(PE_74_io_out_y_im)
  );
  PE PE_75 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_75_clock),
    .io_reset(PE_75_io_reset),
    .io_in_x_re(PE_75_io_in_x_re),
    .io_in_x_im(PE_75_io_in_x_im),
    .io_in_y_re(PE_75_io_in_y_re),
    .io_in_y_im(PE_75_io_in_y_im),
    .io_out_pe_re(PE_75_io_out_pe_re),
    .io_out_pe_im(PE_75_io_out_pe_im),
    .io_out_x_re(PE_75_io_out_x_re),
    .io_out_x_im(PE_75_io_out_x_im),
    .io_out_y_re(PE_75_io_out_y_re),
    .io_out_y_im(PE_75_io_out_y_im)
  );
  PE PE_76 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_76_clock),
    .io_reset(PE_76_io_reset),
    .io_in_x_re(PE_76_io_in_x_re),
    .io_in_x_im(PE_76_io_in_x_im),
    .io_in_y_re(PE_76_io_in_y_re),
    .io_in_y_im(PE_76_io_in_y_im),
    .io_out_pe_re(PE_76_io_out_pe_re),
    .io_out_pe_im(PE_76_io_out_pe_im),
    .io_out_x_re(PE_76_io_out_x_re),
    .io_out_x_im(PE_76_io_out_x_im),
    .io_out_y_re(PE_76_io_out_y_re),
    .io_out_y_im(PE_76_io_out_y_im)
  );
  PE PE_77 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_77_clock),
    .io_reset(PE_77_io_reset),
    .io_in_x_re(PE_77_io_in_x_re),
    .io_in_x_im(PE_77_io_in_x_im),
    .io_in_y_re(PE_77_io_in_y_re),
    .io_in_y_im(PE_77_io_in_y_im),
    .io_out_pe_re(PE_77_io_out_pe_re),
    .io_out_pe_im(PE_77_io_out_pe_im),
    .io_out_x_re(PE_77_io_out_x_re),
    .io_out_x_im(PE_77_io_out_x_im),
    .io_out_y_re(PE_77_io_out_y_re),
    .io_out_y_im(PE_77_io_out_y_im)
  );
  PE PE_78 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_78_clock),
    .io_reset(PE_78_io_reset),
    .io_in_x_re(PE_78_io_in_x_re),
    .io_in_x_im(PE_78_io_in_x_im),
    .io_in_y_re(PE_78_io_in_y_re),
    .io_in_y_im(PE_78_io_in_y_im),
    .io_out_pe_re(PE_78_io_out_pe_re),
    .io_out_pe_im(PE_78_io_out_pe_im),
    .io_out_x_re(PE_78_io_out_x_re),
    .io_out_x_im(PE_78_io_out_x_im),
    .io_out_y_re(PE_78_io_out_y_re),
    .io_out_y_im(PE_78_io_out_y_im)
  );
  PE PE_79 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_79_clock),
    .io_reset(PE_79_io_reset),
    .io_in_x_re(PE_79_io_in_x_re),
    .io_in_x_im(PE_79_io_in_x_im),
    .io_in_y_re(PE_79_io_in_y_re),
    .io_in_y_im(PE_79_io_in_y_im),
    .io_out_pe_re(PE_79_io_out_pe_re),
    .io_out_pe_im(PE_79_io_out_pe_im),
    .io_out_x_re(PE_79_io_out_x_re),
    .io_out_x_im(PE_79_io_out_x_im),
    .io_out_y_re(PE_79_io_out_y_re),
    .io_out_y_im(PE_79_io_out_y_im)
  );
  PE PE_80 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_80_clock),
    .io_reset(PE_80_io_reset),
    .io_in_x_re(PE_80_io_in_x_re),
    .io_in_x_im(PE_80_io_in_x_im),
    .io_in_y_re(PE_80_io_in_y_re),
    .io_in_y_im(PE_80_io_in_y_im),
    .io_out_pe_re(PE_80_io_out_pe_re),
    .io_out_pe_im(PE_80_io_out_pe_im),
    .io_out_x_re(PE_80_io_out_x_re),
    .io_out_x_im(PE_80_io_out_x_im),
    .io_out_y_re(PE_80_io_out_y_re),
    .io_out_y_im(PE_80_io_out_y_im)
  );
  PE PE_81 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_81_clock),
    .io_reset(PE_81_io_reset),
    .io_in_x_re(PE_81_io_in_x_re),
    .io_in_x_im(PE_81_io_in_x_im),
    .io_in_y_re(PE_81_io_in_y_re),
    .io_in_y_im(PE_81_io_in_y_im),
    .io_out_pe_re(PE_81_io_out_pe_re),
    .io_out_pe_im(PE_81_io_out_pe_im),
    .io_out_x_re(PE_81_io_out_x_re),
    .io_out_x_im(PE_81_io_out_x_im),
    .io_out_y_re(PE_81_io_out_y_re),
    .io_out_y_im(PE_81_io_out_y_im)
  );
  PE PE_82 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_82_clock),
    .io_reset(PE_82_io_reset),
    .io_in_x_re(PE_82_io_in_x_re),
    .io_in_x_im(PE_82_io_in_x_im),
    .io_in_y_re(PE_82_io_in_y_re),
    .io_in_y_im(PE_82_io_in_y_im),
    .io_out_pe_re(PE_82_io_out_pe_re),
    .io_out_pe_im(PE_82_io_out_pe_im),
    .io_out_x_re(PE_82_io_out_x_re),
    .io_out_x_im(PE_82_io_out_x_im),
    .io_out_y_re(PE_82_io_out_y_re),
    .io_out_y_im(PE_82_io_out_y_im)
  );
  PE PE_83 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_83_clock),
    .io_reset(PE_83_io_reset),
    .io_in_x_re(PE_83_io_in_x_re),
    .io_in_x_im(PE_83_io_in_x_im),
    .io_in_y_re(PE_83_io_in_y_re),
    .io_in_y_im(PE_83_io_in_y_im),
    .io_out_pe_re(PE_83_io_out_pe_re),
    .io_out_pe_im(PE_83_io_out_pe_im),
    .io_out_x_re(PE_83_io_out_x_re),
    .io_out_x_im(PE_83_io_out_x_im),
    .io_out_y_re(PE_83_io_out_y_re),
    .io_out_y_im(PE_83_io_out_y_im)
  );
  PE PE_84 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_84_clock),
    .io_reset(PE_84_io_reset),
    .io_in_x_re(PE_84_io_in_x_re),
    .io_in_x_im(PE_84_io_in_x_im),
    .io_in_y_re(PE_84_io_in_y_re),
    .io_in_y_im(PE_84_io_in_y_im),
    .io_out_pe_re(PE_84_io_out_pe_re),
    .io_out_pe_im(PE_84_io_out_pe_im),
    .io_out_x_re(PE_84_io_out_x_re),
    .io_out_x_im(PE_84_io_out_x_im),
    .io_out_y_re(PE_84_io_out_y_re),
    .io_out_y_im(PE_84_io_out_y_im)
  );
  PE PE_85 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_85_clock),
    .io_reset(PE_85_io_reset),
    .io_in_x_re(PE_85_io_in_x_re),
    .io_in_x_im(PE_85_io_in_x_im),
    .io_in_y_re(PE_85_io_in_y_re),
    .io_in_y_im(PE_85_io_in_y_im),
    .io_out_pe_re(PE_85_io_out_pe_re),
    .io_out_pe_im(PE_85_io_out_pe_im),
    .io_out_x_re(PE_85_io_out_x_re),
    .io_out_x_im(PE_85_io_out_x_im),
    .io_out_y_re(PE_85_io_out_y_re),
    .io_out_y_im(PE_85_io_out_y_im)
  );
  PE PE_86 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_86_clock),
    .io_reset(PE_86_io_reset),
    .io_in_x_re(PE_86_io_in_x_re),
    .io_in_x_im(PE_86_io_in_x_im),
    .io_in_y_re(PE_86_io_in_y_re),
    .io_in_y_im(PE_86_io_in_y_im),
    .io_out_pe_re(PE_86_io_out_pe_re),
    .io_out_pe_im(PE_86_io_out_pe_im),
    .io_out_x_re(PE_86_io_out_x_re),
    .io_out_x_im(PE_86_io_out_x_im),
    .io_out_y_re(PE_86_io_out_y_re),
    .io_out_y_im(PE_86_io_out_y_im)
  );
  PE PE_87 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_87_clock),
    .io_reset(PE_87_io_reset),
    .io_in_x_re(PE_87_io_in_x_re),
    .io_in_x_im(PE_87_io_in_x_im),
    .io_in_y_re(PE_87_io_in_y_re),
    .io_in_y_im(PE_87_io_in_y_im),
    .io_out_pe_re(PE_87_io_out_pe_re),
    .io_out_pe_im(PE_87_io_out_pe_im),
    .io_out_x_re(PE_87_io_out_x_re),
    .io_out_x_im(PE_87_io_out_x_im),
    .io_out_y_re(PE_87_io_out_y_re),
    .io_out_y_im(PE_87_io_out_y_im)
  );
  PE PE_88 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_88_clock),
    .io_reset(PE_88_io_reset),
    .io_in_x_re(PE_88_io_in_x_re),
    .io_in_x_im(PE_88_io_in_x_im),
    .io_in_y_re(PE_88_io_in_y_re),
    .io_in_y_im(PE_88_io_in_y_im),
    .io_out_pe_re(PE_88_io_out_pe_re),
    .io_out_pe_im(PE_88_io_out_pe_im),
    .io_out_x_re(PE_88_io_out_x_re),
    .io_out_x_im(PE_88_io_out_x_im),
    .io_out_y_re(PE_88_io_out_y_re),
    .io_out_y_im(PE_88_io_out_y_im)
  );
  PE PE_89 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_89_clock),
    .io_reset(PE_89_io_reset),
    .io_in_x_re(PE_89_io_in_x_re),
    .io_in_x_im(PE_89_io_in_x_im),
    .io_in_y_re(PE_89_io_in_y_re),
    .io_in_y_im(PE_89_io_in_y_im),
    .io_out_pe_re(PE_89_io_out_pe_re),
    .io_out_pe_im(PE_89_io_out_pe_im),
    .io_out_x_re(PE_89_io_out_x_re),
    .io_out_x_im(PE_89_io_out_x_im),
    .io_out_y_re(PE_89_io_out_y_re),
    .io_out_y_im(PE_89_io_out_y_im)
  );
  PE PE_90 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_90_clock),
    .io_reset(PE_90_io_reset),
    .io_in_x_re(PE_90_io_in_x_re),
    .io_in_x_im(PE_90_io_in_x_im),
    .io_in_y_re(PE_90_io_in_y_re),
    .io_in_y_im(PE_90_io_in_y_im),
    .io_out_pe_re(PE_90_io_out_pe_re),
    .io_out_pe_im(PE_90_io_out_pe_im),
    .io_out_x_re(PE_90_io_out_x_re),
    .io_out_x_im(PE_90_io_out_x_im),
    .io_out_y_re(PE_90_io_out_y_re),
    .io_out_y_im(PE_90_io_out_y_im)
  );
  PE PE_91 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_91_clock),
    .io_reset(PE_91_io_reset),
    .io_in_x_re(PE_91_io_in_x_re),
    .io_in_x_im(PE_91_io_in_x_im),
    .io_in_y_re(PE_91_io_in_y_re),
    .io_in_y_im(PE_91_io_in_y_im),
    .io_out_pe_re(PE_91_io_out_pe_re),
    .io_out_pe_im(PE_91_io_out_pe_im),
    .io_out_x_re(PE_91_io_out_x_re),
    .io_out_x_im(PE_91_io_out_x_im),
    .io_out_y_re(PE_91_io_out_y_re),
    .io_out_y_im(PE_91_io_out_y_im)
  );
  PE PE_92 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_92_clock),
    .io_reset(PE_92_io_reset),
    .io_in_x_re(PE_92_io_in_x_re),
    .io_in_x_im(PE_92_io_in_x_im),
    .io_in_y_re(PE_92_io_in_y_re),
    .io_in_y_im(PE_92_io_in_y_im),
    .io_out_pe_re(PE_92_io_out_pe_re),
    .io_out_pe_im(PE_92_io_out_pe_im),
    .io_out_x_re(PE_92_io_out_x_re),
    .io_out_x_im(PE_92_io_out_x_im),
    .io_out_y_re(PE_92_io_out_y_re),
    .io_out_y_im(PE_92_io_out_y_im)
  );
  PE PE_93 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_93_clock),
    .io_reset(PE_93_io_reset),
    .io_in_x_re(PE_93_io_in_x_re),
    .io_in_x_im(PE_93_io_in_x_im),
    .io_in_y_re(PE_93_io_in_y_re),
    .io_in_y_im(PE_93_io_in_y_im),
    .io_out_pe_re(PE_93_io_out_pe_re),
    .io_out_pe_im(PE_93_io_out_pe_im),
    .io_out_x_re(PE_93_io_out_x_re),
    .io_out_x_im(PE_93_io_out_x_im),
    .io_out_y_re(PE_93_io_out_y_re),
    .io_out_y_im(PE_93_io_out_y_im)
  );
  PE PE_94 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_94_clock),
    .io_reset(PE_94_io_reset),
    .io_in_x_re(PE_94_io_in_x_re),
    .io_in_x_im(PE_94_io_in_x_im),
    .io_in_y_re(PE_94_io_in_y_re),
    .io_in_y_im(PE_94_io_in_y_im),
    .io_out_pe_re(PE_94_io_out_pe_re),
    .io_out_pe_im(PE_94_io_out_pe_im),
    .io_out_x_re(PE_94_io_out_x_re),
    .io_out_x_im(PE_94_io_out_x_im),
    .io_out_y_re(PE_94_io_out_y_re),
    .io_out_y_im(PE_94_io_out_y_im)
  );
  PE PE_95 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_95_clock),
    .io_reset(PE_95_io_reset),
    .io_in_x_re(PE_95_io_in_x_re),
    .io_in_x_im(PE_95_io_in_x_im),
    .io_in_y_re(PE_95_io_in_y_re),
    .io_in_y_im(PE_95_io_in_y_im),
    .io_out_pe_re(PE_95_io_out_pe_re),
    .io_out_pe_im(PE_95_io_out_pe_im),
    .io_out_x_re(PE_95_io_out_x_re),
    .io_out_x_im(PE_95_io_out_x_im),
    .io_out_y_re(PE_95_io_out_y_re),
    .io_out_y_im(PE_95_io_out_y_im)
  );
  PE PE_96 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_96_clock),
    .io_reset(PE_96_io_reset),
    .io_in_x_re(PE_96_io_in_x_re),
    .io_in_x_im(PE_96_io_in_x_im),
    .io_in_y_re(PE_96_io_in_y_re),
    .io_in_y_im(PE_96_io_in_y_im),
    .io_out_pe_re(PE_96_io_out_pe_re),
    .io_out_pe_im(PE_96_io_out_pe_im),
    .io_out_x_re(PE_96_io_out_x_re),
    .io_out_x_im(PE_96_io_out_x_im),
    .io_out_y_re(PE_96_io_out_y_re),
    .io_out_y_im(PE_96_io_out_y_im)
  );
  PE PE_97 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_97_clock),
    .io_reset(PE_97_io_reset),
    .io_in_x_re(PE_97_io_in_x_re),
    .io_in_x_im(PE_97_io_in_x_im),
    .io_in_y_re(PE_97_io_in_y_re),
    .io_in_y_im(PE_97_io_in_y_im),
    .io_out_pe_re(PE_97_io_out_pe_re),
    .io_out_pe_im(PE_97_io_out_pe_im),
    .io_out_x_re(PE_97_io_out_x_re),
    .io_out_x_im(PE_97_io_out_x_im),
    .io_out_y_re(PE_97_io_out_y_re),
    .io_out_y_im(PE_97_io_out_y_im)
  );
  PE PE_98 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_98_clock),
    .io_reset(PE_98_io_reset),
    .io_in_x_re(PE_98_io_in_x_re),
    .io_in_x_im(PE_98_io_in_x_im),
    .io_in_y_re(PE_98_io_in_y_re),
    .io_in_y_im(PE_98_io_in_y_im),
    .io_out_pe_re(PE_98_io_out_pe_re),
    .io_out_pe_im(PE_98_io_out_pe_im),
    .io_out_x_re(PE_98_io_out_x_re),
    .io_out_x_im(PE_98_io_out_x_im),
    .io_out_y_re(PE_98_io_out_y_re),
    .io_out_y_im(PE_98_io_out_y_im)
  );
  PE PE_99 ( // @[Matrix_Mul_V1.scala 86:35]
    .clock(PE_99_clock),
    .io_reset(PE_99_io_reset),
    .io_in_x_re(PE_99_io_in_x_re),
    .io_in_x_im(PE_99_io_in_x_im),
    .io_in_y_re(PE_99_io_in_y_re),
    .io_in_y_im(PE_99_io_in_y_im),
    .io_out_pe_re(PE_99_io_out_pe_re),
    .io_out_pe_im(PE_99_io_out_pe_im),
    .io_out_x_re(PE_99_io_out_x_re),
    .io_out_x_im(PE_99_io_out_x_im),
    .io_out_y_re(PE_99_io_out_y_re),
    .io_out_y_im(PE_99_io_out_y_im)
  );
  assign io_matrixC_0_re = PE_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_0_im = PE_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_1_re = PE_1_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_1_im = PE_1_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_2_re = PE_2_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_2_im = PE_2_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_3_re = PE_3_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_3_im = PE_3_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_4_re = PE_4_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_4_im = PE_4_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_5_re = PE_5_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_5_im = PE_5_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_6_re = PE_6_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_6_im = PE_6_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_7_re = PE_7_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_7_im = PE_7_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_8_re = PE_8_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_8_im = PE_8_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_9_re = PE_9_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_9_im = PE_9_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_10_re = PE_10_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_10_im = PE_10_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_11_re = PE_11_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_11_im = PE_11_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_12_re = PE_12_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_12_im = PE_12_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_13_re = PE_13_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_13_im = PE_13_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_14_re = PE_14_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_14_im = PE_14_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_15_re = PE_15_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_15_im = PE_15_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_16_re = PE_16_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_16_im = PE_16_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_17_re = PE_17_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_17_im = PE_17_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_18_re = PE_18_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_18_im = PE_18_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_19_re = PE_19_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_19_im = PE_19_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_20_re = PE_20_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_20_im = PE_20_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_21_re = PE_21_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_21_im = PE_21_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_22_re = PE_22_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_22_im = PE_22_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_23_re = PE_23_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_23_im = PE_23_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_24_re = PE_24_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_24_im = PE_24_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_25_re = PE_25_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_25_im = PE_25_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_26_re = PE_26_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_26_im = PE_26_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_27_re = PE_27_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_27_im = PE_27_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_28_re = PE_28_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_28_im = PE_28_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_29_re = PE_29_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_29_im = PE_29_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_30_re = PE_30_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_30_im = PE_30_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_31_re = PE_31_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_31_im = PE_31_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_32_re = PE_32_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_32_im = PE_32_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_33_re = PE_33_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_33_im = PE_33_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_34_re = PE_34_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_34_im = PE_34_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_35_re = PE_35_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_35_im = PE_35_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_36_re = PE_36_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_36_im = PE_36_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_37_re = PE_37_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_37_im = PE_37_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_38_re = PE_38_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_38_im = PE_38_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_39_re = PE_39_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_39_im = PE_39_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_40_re = PE_40_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_40_im = PE_40_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_41_re = PE_41_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_41_im = PE_41_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_42_re = PE_42_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_42_im = PE_42_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_43_re = PE_43_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_43_im = PE_43_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_44_re = PE_44_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_44_im = PE_44_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_45_re = PE_45_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_45_im = PE_45_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_46_re = PE_46_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_46_im = PE_46_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_47_re = PE_47_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_47_im = PE_47_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_48_re = PE_48_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_48_im = PE_48_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_49_re = PE_49_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_49_im = PE_49_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_50_re = PE_50_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_50_im = PE_50_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_51_re = PE_51_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_51_im = PE_51_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_52_re = PE_52_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_52_im = PE_52_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_53_re = PE_53_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_53_im = PE_53_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_54_re = PE_54_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_54_im = PE_54_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_55_re = PE_55_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_55_im = PE_55_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_56_re = PE_56_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_56_im = PE_56_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_57_re = PE_57_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_57_im = PE_57_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_58_re = PE_58_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_58_im = PE_58_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_59_re = PE_59_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_59_im = PE_59_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_60_re = PE_60_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_60_im = PE_60_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_61_re = PE_61_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_61_im = PE_61_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_62_re = PE_62_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_62_im = PE_62_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_63_re = PE_63_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_63_im = PE_63_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_64_re = PE_64_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_64_im = PE_64_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_65_re = PE_65_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_65_im = PE_65_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_66_re = PE_66_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_66_im = PE_66_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_67_re = PE_67_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_67_im = PE_67_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_68_re = PE_68_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_68_im = PE_68_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_69_re = PE_69_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_69_im = PE_69_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_70_re = PE_70_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_70_im = PE_70_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_71_re = PE_71_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_71_im = PE_71_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_72_re = PE_72_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_72_im = PE_72_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_73_re = PE_73_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_73_im = PE_73_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_74_re = PE_74_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_74_im = PE_74_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_75_re = PE_75_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_75_im = PE_75_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_76_re = PE_76_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_76_im = PE_76_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_77_re = PE_77_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_77_im = PE_77_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_78_re = PE_78_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_78_im = PE_78_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_79_re = PE_79_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_79_im = PE_79_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_80_re = PE_80_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_80_im = PE_80_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_81_re = PE_81_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_81_im = PE_81_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_82_re = PE_82_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_82_im = PE_82_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_83_re = PE_83_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_83_im = PE_83_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_84_re = PE_84_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_84_im = PE_84_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_85_re = PE_85_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_85_im = PE_85_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_86_re = PE_86_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_86_im = PE_86_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_87_re = PE_87_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_87_im = PE_87_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_88_re = PE_88_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_88_im = PE_88_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_89_re = PE_89_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_89_im = PE_89_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_90_re = PE_90_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_90_im = PE_90_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_91_re = PE_91_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_91_im = PE_91_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_92_re = PE_92_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_92_im = PE_92_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_93_re = PE_93_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_93_im = PE_93_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_94_re = PE_94_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_94_im = PE_94_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_95_re = PE_95_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_95_im = PE_95_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_96_re = PE_96_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_96_im = PE_96_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_97_re = PE_97_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_97_im = PE_97_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_98_re = PE_98_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_98_im = PE_98_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_99_re = PE_99_io_out_pe_re; // @[Matrix_Mul_V1.scala 195:19]
  assign io_matrixC_99_im = PE_99_io_out_pe_im; // @[Matrix_Mul_V1.scala 195:19]
  assign io_valid = input_point >= 6'h1c; // @[Matrix_Mul_V1.scala 188:20]
  assign PE_clock = clock;
  assign PE_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_io_in_x_re = input_point < 6'h13 ? $signed(_GEN_1183) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_io_in_x_im = input_point < 6'h13 ? $signed(_GEN_993) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_io_in_y_re = _T ? $signed(_GEN_5003) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_io_in_y_im = _T ? $signed(_GEN_4813) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_1_clock = clock;
  assign PE_1_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_1_io_in_x_re = PE_io_out_x_re; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_1_io_in_x_im = PE_io_out_x_im; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_1_io_in_y_re = _T ? $signed(_GEN_5383) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_1_io_in_y_im = _T ? $signed(_GEN_5193) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_2_clock = clock;
  assign PE_2_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_2_io_in_x_re = PE_1_io_out_x_re; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_2_io_in_x_im = PE_1_io_out_x_im; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_2_io_in_y_re = _T ? $signed(_GEN_5763) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_2_io_in_y_im = _T ? $signed(_GEN_5573) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_3_clock = clock;
  assign PE_3_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_3_io_in_x_re = PE_2_io_out_x_re; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_3_io_in_x_im = PE_2_io_out_x_im; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_3_io_in_y_re = _T ? $signed(_GEN_6143) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_3_io_in_y_im = _T ? $signed(_GEN_5953) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_4_clock = clock;
  assign PE_4_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_4_io_in_x_re = PE_3_io_out_x_re; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_4_io_in_x_im = PE_3_io_out_x_im; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_4_io_in_y_re = _T ? $signed(_GEN_6523) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_4_io_in_y_im = _T ? $signed(_GEN_6333) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_5_clock = clock;
  assign PE_5_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_5_io_in_x_re = PE_4_io_out_x_re; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_5_io_in_x_im = PE_4_io_out_x_im; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_5_io_in_y_re = _T ? $signed(_GEN_6903) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_5_io_in_y_im = _T ? $signed(_GEN_6713) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_6_clock = clock;
  assign PE_6_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_6_io_in_x_re = PE_5_io_out_x_re; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_6_io_in_x_im = PE_5_io_out_x_im; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_6_io_in_y_re = _T ? $signed(_GEN_7283) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_6_io_in_y_im = _T ? $signed(_GEN_7093) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_7_clock = clock;
  assign PE_7_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_7_io_in_x_re = PE_6_io_out_x_re; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_7_io_in_x_im = PE_6_io_out_x_im; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_7_io_in_y_re = _T ? $signed(_GEN_7663) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_7_io_in_y_im = _T ? $signed(_GEN_7473) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_8_clock = clock;
  assign PE_8_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_8_io_in_x_re = PE_7_io_out_x_re; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_8_io_in_x_im = PE_7_io_out_x_im; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_8_io_in_y_re = _T ? $signed(_GEN_8043) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_8_io_in_y_im = _T ? $signed(_GEN_7853) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_9_clock = clock;
  assign PE_9_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_9_io_in_x_re = PE_8_io_out_x_re; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_9_io_in_x_im = PE_8_io_out_x_im; // @[Matrix_Mul_V1.scala 178:17]
  assign PE_9_io_in_y_re = _T ? $signed(_GEN_8423) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 167:22]
  assign PE_9_io_in_y_im = _T ? $signed(_GEN_8233) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 159:37 162:19 168:22]
  assign PE_10_clock = clock;
  assign PE_10_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_10_io_in_x_re = input_point < 6'h13 ? $signed(_GEN_1563) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_10_io_in_x_im = input_point < 6'h13 ? $signed(_GEN_1373) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_10_io_in_y_re = PE_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_10_io_in_y_im = PE_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_11_clock = clock;
  assign PE_11_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_11_io_in_x_re = PE_10_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_11_io_in_x_im = PE_10_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_11_io_in_y_re = PE_1_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_11_io_in_y_im = PE_1_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_12_clock = clock;
  assign PE_12_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_12_io_in_x_re = PE_11_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_12_io_in_x_im = PE_11_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_12_io_in_y_re = PE_2_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_12_io_in_y_im = PE_2_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_13_clock = clock;
  assign PE_13_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_13_io_in_x_re = PE_12_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_13_io_in_x_im = PE_12_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_13_io_in_y_re = PE_3_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_13_io_in_y_im = PE_3_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_14_clock = clock;
  assign PE_14_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_14_io_in_x_re = PE_13_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_14_io_in_x_im = PE_13_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_14_io_in_y_re = PE_4_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_14_io_in_y_im = PE_4_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_15_clock = clock;
  assign PE_15_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_15_io_in_x_re = PE_14_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_15_io_in_x_im = PE_14_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_15_io_in_y_re = PE_5_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_15_io_in_y_im = PE_5_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_16_clock = clock;
  assign PE_16_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_16_io_in_x_re = PE_15_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_16_io_in_x_im = PE_15_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_16_io_in_y_re = PE_6_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_16_io_in_y_im = PE_6_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_17_clock = clock;
  assign PE_17_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_17_io_in_x_re = PE_16_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_17_io_in_x_im = PE_16_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_17_io_in_y_re = PE_7_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_17_io_in_y_im = PE_7_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_18_clock = clock;
  assign PE_18_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_18_io_in_x_re = PE_17_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_18_io_in_x_im = PE_17_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_18_io_in_y_re = PE_8_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_18_io_in_y_im = PE_8_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_19_clock = clock;
  assign PE_19_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_19_io_in_x_re = PE_18_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_19_io_in_x_im = PE_18_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_19_io_in_y_re = PE_9_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_19_io_in_y_im = PE_9_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_20_clock = clock;
  assign PE_20_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_20_io_in_x_re = input_point < 6'h13 ? $signed(_GEN_1943) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_20_io_in_x_im = input_point < 6'h13 ? $signed(_GEN_1753) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_20_io_in_y_re = PE_10_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_20_io_in_y_im = PE_10_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_21_clock = clock;
  assign PE_21_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_21_io_in_x_re = PE_20_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_21_io_in_x_im = PE_20_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_21_io_in_y_re = PE_11_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_21_io_in_y_im = PE_11_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_22_clock = clock;
  assign PE_22_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_22_io_in_x_re = PE_21_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_22_io_in_x_im = PE_21_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_22_io_in_y_re = PE_12_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_22_io_in_y_im = PE_12_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_23_clock = clock;
  assign PE_23_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_23_io_in_x_re = PE_22_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_23_io_in_x_im = PE_22_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_23_io_in_y_re = PE_13_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_23_io_in_y_im = PE_13_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_24_clock = clock;
  assign PE_24_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_24_io_in_x_re = PE_23_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_24_io_in_x_im = PE_23_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_24_io_in_y_re = PE_14_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_24_io_in_y_im = PE_14_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_25_clock = clock;
  assign PE_25_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_25_io_in_x_re = PE_24_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_25_io_in_x_im = PE_24_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_25_io_in_y_re = PE_15_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_25_io_in_y_im = PE_15_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_26_clock = clock;
  assign PE_26_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_26_io_in_x_re = PE_25_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_26_io_in_x_im = PE_25_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_26_io_in_y_re = PE_16_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_26_io_in_y_im = PE_16_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_27_clock = clock;
  assign PE_27_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_27_io_in_x_re = PE_26_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_27_io_in_x_im = PE_26_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_27_io_in_y_re = PE_17_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_27_io_in_y_im = PE_17_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_28_clock = clock;
  assign PE_28_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_28_io_in_x_re = PE_27_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_28_io_in_x_im = PE_27_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_28_io_in_y_re = PE_18_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_28_io_in_y_im = PE_18_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_29_clock = clock;
  assign PE_29_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_29_io_in_x_re = PE_28_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_29_io_in_x_im = PE_28_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_29_io_in_y_re = PE_19_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_29_io_in_y_im = PE_19_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_30_clock = clock;
  assign PE_30_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_30_io_in_x_re = input_point < 6'h13 ? $signed(_GEN_2323) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_30_io_in_x_im = input_point < 6'h13 ? $signed(_GEN_2133) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_30_io_in_y_re = PE_20_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_30_io_in_y_im = PE_20_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_31_clock = clock;
  assign PE_31_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_31_io_in_x_re = PE_30_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_31_io_in_x_im = PE_30_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_31_io_in_y_re = PE_21_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_31_io_in_y_im = PE_21_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_32_clock = clock;
  assign PE_32_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_32_io_in_x_re = PE_31_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_32_io_in_x_im = PE_31_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_32_io_in_y_re = PE_22_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_32_io_in_y_im = PE_22_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_33_clock = clock;
  assign PE_33_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_33_io_in_x_re = PE_32_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_33_io_in_x_im = PE_32_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_33_io_in_y_re = PE_23_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_33_io_in_y_im = PE_23_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_34_clock = clock;
  assign PE_34_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_34_io_in_x_re = PE_33_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_34_io_in_x_im = PE_33_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_34_io_in_y_re = PE_24_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_34_io_in_y_im = PE_24_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_35_clock = clock;
  assign PE_35_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_35_io_in_x_re = PE_34_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_35_io_in_x_im = PE_34_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_35_io_in_y_re = PE_25_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_35_io_in_y_im = PE_25_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_36_clock = clock;
  assign PE_36_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_36_io_in_x_re = PE_35_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_36_io_in_x_im = PE_35_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_36_io_in_y_re = PE_26_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_36_io_in_y_im = PE_26_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_37_clock = clock;
  assign PE_37_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_37_io_in_x_re = PE_36_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_37_io_in_x_im = PE_36_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_37_io_in_y_re = PE_27_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_37_io_in_y_im = PE_27_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_38_clock = clock;
  assign PE_38_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_38_io_in_x_re = PE_37_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_38_io_in_x_im = PE_37_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_38_io_in_y_re = PE_28_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_38_io_in_y_im = PE_28_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_39_clock = clock;
  assign PE_39_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_39_io_in_x_re = PE_38_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_39_io_in_x_im = PE_38_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_39_io_in_y_re = PE_29_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_39_io_in_y_im = PE_29_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_40_clock = clock;
  assign PE_40_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_40_io_in_x_re = input_point < 6'h13 ? $signed(_GEN_2703) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_40_io_in_x_im = input_point < 6'h13 ? $signed(_GEN_2513) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_40_io_in_y_re = PE_30_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_40_io_in_y_im = PE_30_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_41_clock = clock;
  assign PE_41_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_41_io_in_x_re = PE_40_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_41_io_in_x_im = PE_40_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_41_io_in_y_re = PE_31_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_41_io_in_y_im = PE_31_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_42_clock = clock;
  assign PE_42_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_42_io_in_x_re = PE_41_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_42_io_in_x_im = PE_41_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_42_io_in_y_re = PE_32_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_42_io_in_y_im = PE_32_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_43_clock = clock;
  assign PE_43_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_43_io_in_x_re = PE_42_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_43_io_in_x_im = PE_42_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_43_io_in_y_re = PE_33_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_43_io_in_y_im = PE_33_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_44_clock = clock;
  assign PE_44_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_44_io_in_x_re = PE_43_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_44_io_in_x_im = PE_43_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_44_io_in_y_re = PE_34_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_44_io_in_y_im = PE_34_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_45_clock = clock;
  assign PE_45_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_45_io_in_x_re = PE_44_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_45_io_in_x_im = PE_44_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_45_io_in_y_re = PE_35_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_45_io_in_y_im = PE_35_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_46_clock = clock;
  assign PE_46_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_46_io_in_x_re = PE_45_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_46_io_in_x_im = PE_45_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_46_io_in_y_re = PE_36_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_46_io_in_y_im = PE_36_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_47_clock = clock;
  assign PE_47_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_47_io_in_x_re = PE_46_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_47_io_in_x_im = PE_46_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_47_io_in_y_re = PE_37_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_47_io_in_y_im = PE_37_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_48_clock = clock;
  assign PE_48_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_48_io_in_x_re = PE_47_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_48_io_in_x_im = PE_47_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_48_io_in_y_re = PE_38_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_48_io_in_y_im = PE_38_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_49_clock = clock;
  assign PE_49_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_49_io_in_x_re = PE_48_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_49_io_in_x_im = PE_48_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_49_io_in_y_re = PE_39_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_49_io_in_y_im = PE_39_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_50_clock = clock;
  assign PE_50_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_50_io_in_x_re = input_point < 6'h13 ? $signed(_GEN_3083) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_50_io_in_x_im = input_point < 6'h13 ? $signed(_GEN_2893) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_50_io_in_y_re = PE_40_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_50_io_in_y_im = PE_40_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_51_clock = clock;
  assign PE_51_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_51_io_in_x_re = PE_50_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_51_io_in_x_im = PE_50_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_51_io_in_y_re = PE_41_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_51_io_in_y_im = PE_41_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_52_clock = clock;
  assign PE_52_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_52_io_in_x_re = PE_51_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_52_io_in_x_im = PE_51_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_52_io_in_y_re = PE_42_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_52_io_in_y_im = PE_42_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_53_clock = clock;
  assign PE_53_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_53_io_in_x_re = PE_52_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_53_io_in_x_im = PE_52_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_53_io_in_y_re = PE_43_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_53_io_in_y_im = PE_43_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_54_clock = clock;
  assign PE_54_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_54_io_in_x_re = PE_53_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_54_io_in_x_im = PE_53_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_54_io_in_y_re = PE_44_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_54_io_in_y_im = PE_44_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_55_clock = clock;
  assign PE_55_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_55_io_in_x_re = PE_54_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_55_io_in_x_im = PE_54_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_55_io_in_y_re = PE_45_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_55_io_in_y_im = PE_45_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_56_clock = clock;
  assign PE_56_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_56_io_in_x_re = PE_55_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_56_io_in_x_im = PE_55_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_56_io_in_y_re = PE_46_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_56_io_in_y_im = PE_46_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_57_clock = clock;
  assign PE_57_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_57_io_in_x_re = PE_56_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_57_io_in_x_im = PE_56_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_57_io_in_y_re = PE_47_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_57_io_in_y_im = PE_47_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_58_clock = clock;
  assign PE_58_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_58_io_in_x_re = PE_57_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_58_io_in_x_im = PE_57_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_58_io_in_y_re = PE_48_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_58_io_in_y_im = PE_48_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_59_clock = clock;
  assign PE_59_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_59_io_in_x_re = PE_58_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_59_io_in_x_im = PE_58_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_59_io_in_y_re = PE_49_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_59_io_in_y_im = PE_49_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_60_clock = clock;
  assign PE_60_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_60_io_in_x_re = input_point < 6'h13 ? $signed(_GEN_3463) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_60_io_in_x_im = input_point < 6'h13 ? $signed(_GEN_3273) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_60_io_in_y_re = PE_50_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_60_io_in_y_im = PE_50_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_61_clock = clock;
  assign PE_61_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_61_io_in_x_re = PE_60_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_61_io_in_x_im = PE_60_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_61_io_in_y_re = PE_51_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_61_io_in_y_im = PE_51_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_62_clock = clock;
  assign PE_62_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_62_io_in_x_re = PE_61_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_62_io_in_x_im = PE_61_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_62_io_in_y_re = PE_52_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_62_io_in_y_im = PE_52_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_63_clock = clock;
  assign PE_63_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_63_io_in_x_re = PE_62_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_63_io_in_x_im = PE_62_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_63_io_in_y_re = PE_53_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_63_io_in_y_im = PE_53_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_64_clock = clock;
  assign PE_64_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_64_io_in_x_re = PE_63_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_64_io_in_x_im = PE_63_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_64_io_in_y_re = PE_54_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_64_io_in_y_im = PE_54_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_65_clock = clock;
  assign PE_65_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_65_io_in_x_re = PE_64_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_65_io_in_x_im = PE_64_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_65_io_in_y_re = PE_55_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_65_io_in_y_im = PE_55_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_66_clock = clock;
  assign PE_66_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_66_io_in_x_re = PE_65_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_66_io_in_x_im = PE_65_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_66_io_in_y_re = PE_56_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_66_io_in_y_im = PE_56_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_67_clock = clock;
  assign PE_67_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_67_io_in_x_re = PE_66_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_67_io_in_x_im = PE_66_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_67_io_in_y_re = PE_57_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_67_io_in_y_im = PE_57_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_68_clock = clock;
  assign PE_68_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_68_io_in_x_re = PE_67_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_68_io_in_x_im = PE_67_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_68_io_in_y_re = PE_58_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_68_io_in_y_im = PE_58_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_69_clock = clock;
  assign PE_69_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_69_io_in_x_re = PE_68_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_69_io_in_x_im = PE_68_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_69_io_in_y_re = PE_59_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_69_io_in_y_im = PE_59_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_70_clock = clock;
  assign PE_70_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_70_io_in_x_re = input_point < 6'h13 ? $signed(_GEN_3843) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_70_io_in_x_im = input_point < 6'h13 ? $signed(_GEN_3653) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_70_io_in_y_re = PE_60_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_70_io_in_y_im = PE_60_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_71_clock = clock;
  assign PE_71_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_71_io_in_x_re = PE_70_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_71_io_in_x_im = PE_70_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_71_io_in_y_re = PE_61_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_71_io_in_y_im = PE_61_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_72_clock = clock;
  assign PE_72_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_72_io_in_x_re = PE_71_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_72_io_in_x_im = PE_71_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_72_io_in_y_re = PE_62_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_72_io_in_y_im = PE_62_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_73_clock = clock;
  assign PE_73_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_73_io_in_x_re = PE_72_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_73_io_in_x_im = PE_72_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_73_io_in_y_re = PE_63_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_73_io_in_y_im = PE_63_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_74_clock = clock;
  assign PE_74_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_74_io_in_x_re = PE_73_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_74_io_in_x_im = PE_73_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_74_io_in_y_re = PE_64_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_74_io_in_y_im = PE_64_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_75_clock = clock;
  assign PE_75_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_75_io_in_x_re = PE_74_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_75_io_in_x_im = PE_74_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_75_io_in_y_re = PE_65_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_75_io_in_y_im = PE_65_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_76_clock = clock;
  assign PE_76_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_76_io_in_x_re = PE_75_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_76_io_in_x_im = PE_75_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_76_io_in_y_re = PE_66_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_76_io_in_y_im = PE_66_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_77_clock = clock;
  assign PE_77_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_77_io_in_x_re = PE_76_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_77_io_in_x_im = PE_76_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_77_io_in_y_re = PE_67_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_77_io_in_y_im = PE_67_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_78_clock = clock;
  assign PE_78_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_78_io_in_x_re = PE_77_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_78_io_in_x_im = PE_77_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_78_io_in_y_re = PE_68_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_78_io_in_y_im = PE_68_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_79_clock = clock;
  assign PE_79_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_79_io_in_x_re = PE_78_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_79_io_in_x_im = PE_78_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_79_io_in_y_re = PE_69_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_79_io_in_y_im = PE_69_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_80_clock = clock;
  assign PE_80_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_80_io_in_x_re = input_point < 6'h13 ? $signed(_GEN_4223) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_80_io_in_x_im = input_point < 6'h13 ? $signed(_GEN_4033) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_80_io_in_y_re = PE_70_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_80_io_in_y_im = PE_70_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_81_clock = clock;
  assign PE_81_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_81_io_in_x_re = PE_80_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_81_io_in_x_im = PE_80_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_81_io_in_y_re = PE_71_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_81_io_in_y_im = PE_71_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_82_clock = clock;
  assign PE_82_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_82_io_in_x_re = PE_81_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_82_io_in_x_im = PE_81_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_82_io_in_y_re = PE_72_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_82_io_in_y_im = PE_72_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_83_clock = clock;
  assign PE_83_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_83_io_in_x_re = PE_82_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_83_io_in_x_im = PE_82_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_83_io_in_y_re = PE_73_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_83_io_in_y_im = PE_73_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_84_clock = clock;
  assign PE_84_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_84_io_in_x_re = PE_83_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_84_io_in_x_im = PE_83_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_84_io_in_y_re = PE_74_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_84_io_in_y_im = PE_74_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_85_clock = clock;
  assign PE_85_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_85_io_in_x_re = PE_84_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_85_io_in_x_im = PE_84_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_85_io_in_y_re = PE_75_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_85_io_in_y_im = PE_75_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_86_clock = clock;
  assign PE_86_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_86_io_in_x_re = PE_85_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_86_io_in_x_im = PE_85_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_86_io_in_y_re = PE_76_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_86_io_in_y_im = PE_76_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_87_clock = clock;
  assign PE_87_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_87_io_in_x_re = PE_86_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_87_io_in_x_im = PE_86_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_87_io_in_y_re = PE_77_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_87_io_in_y_im = PE_77_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_88_clock = clock;
  assign PE_88_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_88_io_in_x_re = PE_87_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_88_io_in_x_im = PE_87_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_88_io_in_y_re = PE_78_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_88_io_in_y_im = PE_78_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_89_clock = clock;
  assign PE_89_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_89_io_in_x_re = PE_88_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_89_io_in_x_im = PE_88_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_89_io_in_y_re = PE_79_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_89_io_in_y_im = PE_79_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_90_clock = clock;
  assign PE_90_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_90_io_in_x_re = input_point < 6'h13 ? $signed(_GEN_4603) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 153:30]
  assign PE_90_io_in_x_im = input_point < 6'h13 ? $signed(_GEN_4413) : $signed(32'sh0); // @[Matrix_Mul_V1.scala 145:37 148:27 154:30]
  assign PE_90_io_in_y_re = PE_80_io_out_y_re; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_90_io_in_y_im = PE_80_io_out_y_im; // @[Matrix_Mul_V1.scala 175:25]
  assign PE_91_clock = clock;
  assign PE_91_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_91_io_in_x_re = PE_90_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_91_io_in_x_im = PE_90_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_91_io_in_y_re = PE_81_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_91_io_in_y_im = PE_81_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_92_clock = clock;
  assign PE_92_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_92_io_in_x_re = PE_91_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_92_io_in_x_im = PE_91_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_92_io_in_y_re = PE_82_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_92_io_in_y_im = PE_82_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_93_clock = clock;
  assign PE_93_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_93_io_in_x_re = PE_92_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_93_io_in_x_im = PE_92_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_93_io_in_y_re = PE_83_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_93_io_in_y_im = PE_83_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_94_clock = clock;
  assign PE_94_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_94_io_in_x_re = PE_93_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_94_io_in_x_im = PE_93_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_94_io_in_y_re = PE_84_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_94_io_in_y_im = PE_84_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_95_clock = clock;
  assign PE_95_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_95_io_in_x_re = PE_94_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_95_io_in_x_im = PE_94_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_95_io_in_y_re = PE_85_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_95_io_in_y_im = PE_85_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_96_clock = clock;
  assign PE_96_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_96_io_in_x_re = PE_95_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_96_io_in_x_im = PE_95_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_96_io_in_y_re = PE_86_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_96_io_in_y_im = PE_86_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_97_clock = clock;
  assign PE_97_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_97_io_in_x_re = PE_96_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_97_io_in_x_im = PE_96_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_97_io_in_y_re = PE_87_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_97_io_in_y_im = PE_87_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_98_clock = clock;
  assign PE_98_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_98_io_in_x_re = PE_97_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_98_io_in_x_im = PE_97_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_98_io_in_y_re = PE_88_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_98_io_in_y_im = PE_88_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_99_clock = clock;
  assign PE_99_io_reset = io_reset | io_ready; // @[Matrix_Mul_V1.scala 89:18 101:20]
  assign PE_99_io_in_x_re = PE_98_io_out_x_re; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_99_io_in_x_im = PE_98_io_out_x_im; // @[Matrix_Mul_V1.scala 183:27]
  assign PE_99_io_in_y_re = PE_89_io_out_y_re; // @[Matrix_Mul_V1.scala 182:27]
  assign PE_99_io_in_y_im = PE_89_io_out_y_im; // @[Matrix_Mul_V1.scala 182:27]
  always @(posedge clock) begin
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_0_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_0_re <= io_matrixA_0_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_0_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_0_im <= io_matrixA_0_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_1_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_1_re <= io_matrixA_1_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_1_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_1_im <= io_matrixA_1_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_2_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_2_re <= io_matrixA_2_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_2_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_2_im <= io_matrixA_2_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_3_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_3_re <= io_matrixA_3_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_3_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_3_im <= io_matrixA_3_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_4_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_4_re <= io_matrixA_4_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_4_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_4_im <= io_matrixA_4_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_5_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_5_re <= io_matrixA_5_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_5_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_5_im <= io_matrixA_5_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_6_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_6_re <= io_matrixA_6_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_6_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_6_im <= io_matrixA_6_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_7_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_7_re <= io_matrixA_7_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_7_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_7_im <= io_matrixA_7_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_8_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_8_re <= io_matrixA_8_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_8_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_8_im <= io_matrixA_8_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_9_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_9_re <= io_matrixA_9_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_9_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_9_im <= io_matrixA_9_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_10_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_10_re <= io_matrixA_10_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_10_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_10_im <= io_matrixA_10_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_11_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_11_re <= io_matrixA_11_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_11_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_11_im <= io_matrixA_11_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_12_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_12_re <= io_matrixA_12_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_12_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_12_im <= io_matrixA_12_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_13_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_13_re <= io_matrixA_13_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_13_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_13_im <= io_matrixA_13_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_14_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_14_re <= io_matrixA_14_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_14_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_14_im <= io_matrixA_14_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_15_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_15_re <= io_matrixA_15_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_15_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_15_im <= io_matrixA_15_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_16_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_16_re <= io_matrixA_16_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_16_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_16_im <= io_matrixA_16_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_17_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_17_re <= io_matrixA_17_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_17_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_17_im <= io_matrixA_17_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_18_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_18_re <= io_matrixA_18_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_18_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_18_im <= io_matrixA_18_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_19_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_19_re <= io_matrixA_19_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_19_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_19_im <= io_matrixA_19_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_20_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_20_re <= io_matrixA_20_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_20_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_20_im <= io_matrixA_20_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_21_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_21_re <= io_matrixA_21_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_21_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_21_im <= io_matrixA_21_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_22_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_22_re <= io_matrixA_22_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_22_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_22_im <= io_matrixA_22_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_23_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_23_re <= io_matrixA_23_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_23_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_23_im <= io_matrixA_23_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_24_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_24_re <= io_matrixA_24_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_24_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_24_im <= io_matrixA_24_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_25_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_25_re <= io_matrixA_25_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_25_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_25_im <= io_matrixA_25_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_26_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_26_re <= io_matrixA_26_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_26_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_26_im <= io_matrixA_26_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_27_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_27_re <= io_matrixA_27_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_27_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_27_im <= io_matrixA_27_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_28_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_28_re <= io_matrixA_28_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_28_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_28_im <= io_matrixA_28_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_29_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_29_re <= io_matrixA_29_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_29_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_29_im <= io_matrixA_29_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_30_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_30_re <= io_matrixA_30_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_30_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_30_im <= io_matrixA_30_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_31_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_31_re <= io_matrixA_31_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_31_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_31_im <= io_matrixA_31_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_32_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_32_re <= io_matrixA_32_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_32_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_32_im <= io_matrixA_32_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_33_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_33_re <= io_matrixA_33_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_33_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_33_im <= io_matrixA_33_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_34_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_34_re <= io_matrixA_34_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_34_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_34_im <= io_matrixA_34_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_35_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_35_re <= io_matrixA_35_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_35_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_35_im <= io_matrixA_35_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_36_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_36_re <= io_matrixA_36_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_36_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_36_im <= io_matrixA_36_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_37_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_37_re <= io_matrixA_37_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_37_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_37_im <= io_matrixA_37_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_38_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_38_re <= io_matrixA_38_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_38_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_38_im <= io_matrixA_38_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_39_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_39_re <= io_matrixA_39_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_39_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_39_im <= io_matrixA_39_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_40_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_40_re <= io_matrixA_40_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_40_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_40_im <= io_matrixA_40_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_41_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_41_re <= io_matrixA_41_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_41_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_41_im <= io_matrixA_41_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_42_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_42_re <= io_matrixA_42_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_42_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_42_im <= io_matrixA_42_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_43_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_43_re <= io_matrixA_43_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_43_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_43_im <= io_matrixA_43_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_44_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_44_re <= io_matrixA_44_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_44_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_44_im <= io_matrixA_44_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_45_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_45_re <= io_matrixA_45_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_45_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_45_im <= io_matrixA_45_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_46_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_46_re <= io_matrixA_46_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_46_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_46_im <= io_matrixA_46_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_47_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_47_re <= io_matrixA_47_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_47_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_47_im <= io_matrixA_47_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_48_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_48_re <= io_matrixA_48_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_48_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_48_im <= io_matrixA_48_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_49_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_49_re <= io_matrixA_49_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_49_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_49_im <= io_matrixA_49_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_50_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_50_re <= io_matrixA_50_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_50_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_50_im <= io_matrixA_50_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_51_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_51_re <= io_matrixA_51_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_51_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_51_im <= io_matrixA_51_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_52_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_52_re <= io_matrixA_52_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_52_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_52_im <= io_matrixA_52_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_53_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_53_re <= io_matrixA_53_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_53_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_53_im <= io_matrixA_53_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_54_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_54_re <= io_matrixA_54_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_54_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_54_im <= io_matrixA_54_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_55_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_55_re <= io_matrixA_55_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_55_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_55_im <= io_matrixA_55_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_56_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_56_re <= io_matrixA_56_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_56_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_56_im <= io_matrixA_56_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_57_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_57_re <= io_matrixA_57_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_57_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_57_im <= io_matrixA_57_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_58_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_58_re <= io_matrixA_58_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_58_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_58_im <= io_matrixA_58_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_59_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_59_re <= io_matrixA_59_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_59_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_59_im <= io_matrixA_59_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_60_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_60_re <= io_matrixA_60_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_60_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_60_im <= io_matrixA_60_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_61_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_61_re <= io_matrixA_61_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_61_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_61_im <= io_matrixA_61_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_62_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_62_re <= io_matrixA_62_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_62_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_62_im <= io_matrixA_62_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_63_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_63_re <= io_matrixA_63_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_63_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_63_im <= io_matrixA_63_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_64_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_64_re <= io_matrixA_64_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_64_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_64_im <= io_matrixA_64_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_65_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_65_re <= io_matrixA_65_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_65_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_65_im <= io_matrixA_65_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_66_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_66_re <= io_matrixA_66_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_66_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_66_im <= io_matrixA_66_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_67_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_67_re <= io_matrixA_67_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_67_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_67_im <= io_matrixA_67_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_68_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_68_re <= io_matrixA_68_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_68_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_68_im <= io_matrixA_68_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_69_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_69_re <= io_matrixA_69_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_69_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_69_im <= io_matrixA_69_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_70_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_70_re <= io_matrixA_70_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_70_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_70_im <= io_matrixA_70_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_71_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_71_re <= io_matrixA_71_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_71_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_71_im <= io_matrixA_71_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_72_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_72_re <= io_matrixA_72_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_72_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_72_im <= io_matrixA_72_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_73_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_73_re <= io_matrixA_73_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_73_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_73_im <= io_matrixA_73_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_74_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_74_re <= io_matrixA_74_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_74_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_74_im <= io_matrixA_74_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_75_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_75_re <= io_matrixA_75_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_75_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_75_im <= io_matrixA_75_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_76_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_76_re <= io_matrixA_76_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_76_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_76_im <= io_matrixA_76_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_77_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_77_re <= io_matrixA_77_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_77_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_77_im <= io_matrixA_77_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_78_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_78_re <= io_matrixA_78_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_78_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_78_im <= io_matrixA_78_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_79_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_79_re <= io_matrixA_79_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_79_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_79_im <= io_matrixA_79_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_80_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_80_re <= io_matrixA_80_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_80_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_80_im <= io_matrixA_80_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_81_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_81_re <= io_matrixA_81_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_81_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_81_im <= io_matrixA_81_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_82_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_82_re <= io_matrixA_82_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_82_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_82_im <= io_matrixA_82_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_83_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_83_re <= io_matrixA_83_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_83_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_83_im <= io_matrixA_83_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_84_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_84_re <= io_matrixA_84_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_84_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_84_im <= io_matrixA_84_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_85_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_85_re <= io_matrixA_85_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_85_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_85_im <= io_matrixA_85_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_86_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_86_re <= io_matrixA_86_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_86_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_86_im <= io_matrixA_86_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_87_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_87_re <= io_matrixA_87_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_87_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_87_im <= io_matrixA_87_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_88_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_88_re <= io_matrixA_88_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_88_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_88_im <= io_matrixA_88_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_89_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_89_re <= io_matrixA_89_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_89_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_89_im <= io_matrixA_89_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_90_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_90_re <= io_matrixA_90_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_90_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_90_im <= io_matrixA_90_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_91_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_91_re <= io_matrixA_91_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_91_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_91_im <= io_matrixA_91_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_92_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_92_re <= io_matrixA_92_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_92_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_92_im <= io_matrixA_92_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_93_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_93_re <= io_matrixA_93_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_93_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_93_im <= io_matrixA_93_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_94_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_94_re <= io_matrixA_94_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_94_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_94_im <= io_matrixA_94_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_95_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_95_re <= io_matrixA_95_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_95_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_95_im <= io_matrixA_95_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_96_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_96_re <= io_matrixA_96_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_96_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_96_im <= io_matrixA_96_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_97_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_97_re <= io_matrixA_97_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_97_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_97_im <= io_matrixA_97_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_98_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_98_re <= io_matrixA_98_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_98_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_98_im <= io_matrixA_98_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_99_re <= 32'sh0; // @[Matrix_Mul_V1.scala 92:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_99_re <= io_matrixA_99_re; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsA_99_im <= 32'sh0; // @[Matrix_Mul_V1.scala 93:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsA_99_im <= io_matrixA_99_im; // @[Matrix_Mul_V1.scala 105:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_0_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_0_re <= io_matrixB_0_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_0_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_0_im <= io_matrixB_0_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_1_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_1_re <= io_matrixB_1_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_1_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_1_im <= io_matrixB_1_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_2_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_2_re <= io_matrixB_2_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_2_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_2_im <= io_matrixB_2_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_3_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_3_re <= io_matrixB_3_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_3_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_3_im <= io_matrixB_3_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_4_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_4_re <= io_matrixB_4_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_4_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_4_im <= io_matrixB_4_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_5_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_5_re <= io_matrixB_5_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_5_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_5_im <= io_matrixB_5_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_6_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_6_re <= io_matrixB_6_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_6_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_6_im <= io_matrixB_6_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_7_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_7_re <= io_matrixB_7_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_7_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_7_im <= io_matrixB_7_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_8_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_8_re <= io_matrixB_8_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_8_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_8_im <= io_matrixB_8_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_9_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_9_re <= io_matrixB_9_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_9_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_9_im <= io_matrixB_9_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_10_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_10_re <= io_matrixB_10_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_10_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_10_im <= io_matrixB_10_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_11_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_11_re <= io_matrixB_11_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_11_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_11_im <= io_matrixB_11_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_12_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_12_re <= io_matrixB_12_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_12_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_12_im <= io_matrixB_12_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_13_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_13_re <= io_matrixB_13_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_13_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_13_im <= io_matrixB_13_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_14_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_14_re <= io_matrixB_14_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_14_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_14_im <= io_matrixB_14_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_15_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_15_re <= io_matrixB_15_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_15_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_15_im <= io_matrixB_15_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_16_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_16_re <= io_matrixB_16_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_16_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_16_im <= io_matrixB_16_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_17_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_17_re <= io_matrixB_17_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_17_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_17_im <= io_matrixB_17_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_18_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_18_re <= io_matrixB_18_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_18_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_18_im <= io_matrixB_18_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_19_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_19_re <= io_matrixB_19_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_19_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_19_im <= io_matrixB_19_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_20_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_20_re <= io_matrixB_20_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_20_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_20_im <= io_matrixB_20_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_21_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_21_re <= io_matrixB_21_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_21_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_21_im <= io_matrixB_21_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_22_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_22_re <= io_matrixB_22_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_22_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_22_im <= io_matrixB_22_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_23_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_23_re <= io_matrixB_23_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_23_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_23_im <= io_matrixB_23_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_24_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_24_re <= io_matrixB_24_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_24_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_24_im <= io_matrixB_24_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_25_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_25_re <= io_matrixB_25_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_25_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_25_im <= io_matrixB_25_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_26_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_26_re <= io_matrixB_26_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_26_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_26_im <= io_matrixB_26_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_27_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_27_re <= io_matrixB_27_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_27_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_27_im <= io_matrixB_27_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_28_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_28_re <= io_matrixB_28_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_28_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_28_im <= io_matrixB_28_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_29_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_29_re <= io_matrixB_29_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_29_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_29_im <= io_matrixB_29_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_30_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_30_re <= io_matrixB_30_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_30_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_30_im <= io_matrixB_30_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_31_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_31_re <= io_matrixB_31_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_31_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_31_im <= io_matrixB_31_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_32_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_32_re <= io_matrixB_32_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_32_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_32_im <= io_matrixB_32_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_33_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_33_re <= io_matrixB_33_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_33_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_33_im <= io_matrixB_33_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_34_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_34_re <= io_matrixB_34_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_34_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_34_im <= io_matrixB_34_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_35_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_35_re <= io_matrixB_35_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_35_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_35_im <= io_matrixB_35_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_36_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_36_re <= io_matrixB_36_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_36_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_36_im <= io_matrixB_36_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_37_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_37_re <= io_matrixB_37_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_37_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_37_im <= io_matrixB_37_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_38_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_38_re <= io_matrixB_38_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_38_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_38_im <= io_matrixB_38_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_39_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_39_re <= io_matrixB_39_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_39_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_39_im <= io_matrixB_39_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_40_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_40_re <= io_matrixB_40_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_40_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_40_im <= io_matrixB_40_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_41_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_41_re <= io_matrixB_41_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_41_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_41_im <= io_matrixB_41_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_42_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_42_re <= io_matrixB_42_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_42_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_42_im <= io_matrixB_42_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_43_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_43_re <= io_matrixB_43_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_43_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_43_im <= io_matrixB_43_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_44_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_44_re <= io_matrixB_44_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_44_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_44_im <= io_matrixB_44_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_45_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_45_re <= io_matrixB_45_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_45_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_45_im <= io_matrixB_45_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_46_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_46_re <= io_matrixB_46_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_46_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_46_im <= io_matrixB_46_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_47_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_47_re <= io_matrixB_47_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_47_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_47_im <= io_matrixB_47_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_48_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_48_re <= io_matrixB_48_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_48_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_48_im <= io_matrixB_48_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_49_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_49_re <= io_matrixB_49_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_49_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_49_im <= io_matrixB_49_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_50_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_50_re <= io_matrixB_50_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_50_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_50_im <= io_matrixB_50_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_51_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_51_re <= io_matrixB_51_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_51_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_51_im <= io_matrixB_51_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_52_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_52_re <= io_matrixB_52_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_52_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_52_im <= io_matrixB_52_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_53_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_53_re <= io_matrixB_53_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_53_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_53_im <= io_matrixB_53_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_54_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_54_re <= io_matrixB_54_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_54_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_54_im <= io_matrixB_54_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_55_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_55_re <= io_matrixB_55_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_55_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_55_im <= io_matrixB_55_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_56_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_56_re <= io_matrixB_56_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_56_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_56_im <= io_matrixB_56_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_57_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_57_re <= io_matrixB_57_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_57_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_57_im <= io_matrixB_57_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_58_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_58_re <= io_matrixB_58_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_58_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_58_im <= io_matrixB_58_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_59_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_59_re <= io_matrixB_59_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_59_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_59_im <= io_matrixB_59_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_60_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_60_re <= io_matrixB_60_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_60_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_60_im <= io_matrixB_60_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_61_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_61_re <= io_matrixB_61_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_61_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_61_im <= io_matrixB_61_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_62_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_62_re <= io_matrixB_62_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_62_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_62_im <= io_matrixB_62_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_63_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_63_re <= io_matrixB_63_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_63_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_63_im <= io_matrixB_63_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_64_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_64_re <= io_matrixB_64_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_64_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_64_im <= io_matrixB_64_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_65_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_65_re <= io_matrixB_65_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_65_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_65_im <= io_matrixB_65_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_66_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_66_re <= io_matrixB_66_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_66_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_66_im <= io_matrixB_66_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_67_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_67_re <= io_matrixB_67_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_67_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_67_im <= io_matrixB_67_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_68_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_68_re <= io_matrixB_68_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_68_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_68_im <= io_matrixB_68_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_69_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_69_re <= io_matrixB_69_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_69_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_69_im <= io_matrixB_69_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_70_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_70_re <= io_matrixB_70_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_70_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_70_im <= io_matrixB_70_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_71_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_71_re <= io_matrixB_71_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_71_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_71_im <= io_matrixB_71_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_72_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_72_re <= io_matrixB_72_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_72_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_72_im <= io_matrixB_72_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_73_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_73_re <= io_matrixB_73_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_73_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_73_im <= io_matrixB_73_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_74_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_74_re <= io_matrixB_74_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_74_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_74_im <= io_matrixB_74_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_75_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_75_re <= io_matrixB_75_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_75_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_75_im <= io_matrixB_75_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_76_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_76_re <= io_matrixB_76_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_76_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_76_im <= io_matrixB_76_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_77_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_77_re <= io_matrixB_77_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_77_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_77_im <= io_matrixB_77_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_78_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_78_re <= io_matrixB_78_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_78_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_78_im <= io_matrixB_78_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_79_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_79_re <= io_matrixB_79_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_79_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_79_im <= io_matrixB_79_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_80_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_80_re <= io_matrixB_80_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_80_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_80_im <= io_matrixB_80_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_81_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_81_re <= io_matrixB_81_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_81_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_81_im <= io_matrixB_81_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_82_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_82_re <= io_matrixB_82_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_82_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_82_im <= io_matrixB_82_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_83_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_83_re <= io_matrixB_83_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_83_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_83_im <= io_matrixB_83_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_84_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_84_re <= io_matrixB_84_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_84_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_84_im <= io_matrixB_84_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_85_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_85_re <= io_matrixB_85_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_85_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_85_im <= io_matrixB_85_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_86_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_86_re <= io_matrixB_86_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_86_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_86_im <= io_matrixB_86_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_87_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_87_re <= io_matrixB_87_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_87_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_87_im <= io_matrixB_87_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_88_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_88_re <= io_matrixB_88_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_88_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_88_im <= io_matrixB_88_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_89_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_89_re <= io_matrixB_89_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_89_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_89_im <= io_matrixB_89_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_90_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_90_re <= io_matrixB_90_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_90_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_90_im <= io_matrixB_90_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_91_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_91_re <= io_matrixB_91_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_91_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_91_im <= io_matrixB_91_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_92_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_92_re <= io_matrixB_92_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_92_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_92_im <= io_matrixB_92_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_93_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_93_re <= io_matrixB_93_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_93_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_93_im <= io_matrixB_93_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_94_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_94_re <= io_matrixB_94_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_94_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_94_im <= io_matrixB_94_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_95_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_95_re <= io_matrixB_95_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_95_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_95_im <= io_matrixB_95_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_96_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_96_re <= io_matrixB_96_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_96_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_96_im <= io_matrixB_96_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_97_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_97_re <= io_matrixB_97_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_97_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_97_im <= io_matrixB_97_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_98_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_98_re <= io_matrixB_98_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_98_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_98_im <= io_matrixB_98_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_99_re <= 32'sh0; // @[Matrix_Mul_V1.scala 96:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_99_re <= io_matrixB_99_re; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      regsB_99_im <= 32'sh0; // @[Matrix_Mul_V1.scala 97:19]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      regsB_99_im <= io_matrixB_99_im; // @[Matrix_Mul_V1.scala 106:11]
    end
    if (io_reset) begin // @[Matrix_Mul_V1.scala 89:18]
      input_point <= 6'h0; // @[Matrix_Mul_V1.scala 99:17]
    end else if (io_ready) begin // @[Matrix_Mul_V1.scala 103:24]
      input_point <= 6'h0; // @[Matrix_Mul_V1.scala 108:17]
    end else begin
      input_point <= _input_point_T_1; // @[Matrix_Mul_V1.scala 116:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regsA_0_re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regsA_0_im = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regsA_1_re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regsA_1_im = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regsA_2_re = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regsA_2_im = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regsA_3_re = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regsA_3_im = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regsA_4_re = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regsA_4_im = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regsA_5_re = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regsA_5_im = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regsA_6_re = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regsA_6_im = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regsA_7_re = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regsA_7_im = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regsA_8_re = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  regsA_8_im = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regsA_9_re = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  regsA_9_im = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regsA_10_re = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  regsA_10_im = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  regsA_11_re = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  regsA_11_im = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  regsA_12_re = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  regsA_12_im = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  regsA_13_re = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  regsA_13_im = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regsA_14_re = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  regsA_14_im = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regsA_15_re = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  regsA_15_im = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  regsA_16_re = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  regsA_16_im = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  regsA_17_re = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  regsA_17_im = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  regsA_18_re = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  regsA_18_im = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  regsA_19_re = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  regsA_19_im = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  regsA_20_re = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  regsA_20_im = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  regsA_21_re = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  regsA_21_im = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  regsA_22_re = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  regsA_22_im = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  regsA_23_re = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  regsA_23_im = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  regsA_24_re = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  regsA_24_im = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  regsA_25_re = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  regsA_25_im = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  regsA_26_re = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  regsA_26_im = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  regsA_27_re = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  regsA_27_im = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  regsA_28_re = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  regsA_28_im = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  regsA_29_re = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  regsA_29_im = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  regsA_30_re = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  regsA_30_im = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  regsA_31_re = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  regsA_31_im = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  regsA_32_re = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  regsA_32_im = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  regsA_33_re = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  regsA_33_im = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  regsA_34_re = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  regsA_34_im = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  regsA_35_re = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  regsA_35_im = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  regsA_36_re = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  regsA_36_im = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  regsA_37_re = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  regsA_37_im = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  regsA_38_re = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  regsA_38_im = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  regsA_39_re = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  regsA_39_im = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  regsA_40_re = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  regsA_40_im = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  regsA_41_re = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  regsA_41_im = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  regsA_42_re = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  regsA_42_im = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  regsA_43_re = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  regsA_43_im = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  regsA_44_re = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  regsA_44_im = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  regsA_45_re = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  regsA_45_im = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  regsA_46_re = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  regsA_46_im = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  regsA_47_re = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  regsA_47_im = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  regsA_48_re = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  regsA_48_im = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  regsA_49_re = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  regsA_49_im = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  regsA_50_re = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  regsA_50_im = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  regsA_51_re = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  regsA_51_im = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  regsA_52_re = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  regsA_52_im = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  regsA_53_re = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  regsA_53_im = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  regsA_54_re = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  regsA_54_im = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  regsA_55_re = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  regsA_55_im = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  regsA_56_re = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  regsA_56_im = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  regsA_57_re = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  regsA_57_im = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  regsA_58_re = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  regsA_58_im = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  regsA_59_re = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  regsA_59_im = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  regsA_60_re = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  regsA_60_im = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  regsA_61_re = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  regsA_61_im = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  regsA_62_re = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  regsA_62_im = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  regsA_63_re = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  regsA_63_im = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  regsA_64_re = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  regsA_64_im = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  regsA_65_re = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  regsA_65_im = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  regsA_66_re = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  regsA_66_im = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  regsA_67_re = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  regsA_67_im = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  regsA_68_re = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  regsA_68_im = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  regsA_69_re = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  regsA_69_im = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  regsA_70_re = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  regsA_70_im = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  regsA_71_re = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  regsA_71_im = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  regsA_72_re = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  regsA_72_im = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  regsA_73_re = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  regsA_73_im = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  regsA_74_re = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  regsA_74_im = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  regsA_75_re = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  regsA_75_im = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  regsA_76_re = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  regsA_76_im = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  regsA_77_re = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  regsA_77_im = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  regsA_78_re = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  regsA_78_im = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  regsA_79_re = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  regsA_79_im = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  regsA_80_re = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  regsA_80_im = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  regsA_81_re = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  regsA_81_im = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  regsA_82_re = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  regsA_82_im = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  regsA_83_re = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  regsA_83_im = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  regsA_84_re = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  regsA_84_im = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  regsA_85_re = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  regsA_85_im = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  regsA_86_re = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  regsA_86_im = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  regsA_87_re = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  regsA_87_im = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  regsA_88_re = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  regsA_88_im = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  regsA_89_re = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  regsA_89_im = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  regsA_90_re = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  regsA_90_im = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  regsA_91_re = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  regsA_91_im = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  regsA_92_re = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  regsA_92_im = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  regsA_93_re = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  regsA_93_im = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  regsA_94_re = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  regsA_94_im = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  regsA_95_re = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  regsA_95_im = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  regsA_96_re = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  regsA_96_im = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  regsA_97_re = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  regsA_97_im = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  regsA_98_re = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  regsA_98_im = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  regsA_99_re = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  regsA_99_im = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  regsB_0_re = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  regsB_0_im = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  regsB_1_re = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  regsB_1_im = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  regsB_2_re = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  regsB_2_im = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  regsB_3_re = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  regsB_3_im = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  regsB_4_re = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  regsB_4_im = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  regsB_5_re = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  regsB_5_im = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  regsB_6_re = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  regsB_6_im = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  regsB_7_re = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  regsB_7_im = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  regsB_8_re = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  regsB_8_im = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  regsB_9_re = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  regsB_9_im = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  regsB_10_re = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  regsB_10_im = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  regsB_11_re = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  regsB_11_im = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  regsB_12_re = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  regsB_12_im = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  regsB_13_re = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  regsB_13_im = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  regsB_14_re = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  regsB_14_im = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  regsB_15_re = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  regsB_15_im = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  regsB_16_re = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  regsB_16_im = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  regsB_17_re = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  regsB_17_im = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  regsB_18_re = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  regsB_18_im = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  regsB_19_re = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  regsB_19_im = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  regsB_20_re = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  regsB_20_im = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  regsB_21_re = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  regsB_21_im = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  regsB_22_re = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  regsB_22_im = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  regsB_23_re = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  regsB_23_im = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  regsB_24_re = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  regsB_24_im = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  regsB_25_re = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  regsB_25_im = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  regsB_26_re = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  regsB_26_im = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  regsB_27_re = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  regsB_27_im = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  regsB_28_re = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  regsB_28_im = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  regsB_29_re = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  regsB_29_im = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  regsB_30_re = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  regsB_30_im = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  regsB_31_re = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  regsB_31_im = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  regsB_32_re = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  regsB_32_im = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  regsB_33_re = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  regsB_33_im = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  regsB_34_re = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  regsB_34_im = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  regsB_35_re = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  regsB_35_im = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  regsB_36_re = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  regsB_36_im = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  regsB_37_re = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  regsB_37_im = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  regsB_38_re = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  regsB_38_im = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  regsB_39_re = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  regsB_39_im = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  regsB_40_re = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  regsB_40_im = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  regsB_41_re = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  regsB_41_im = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  regsB_42_re = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  regsB_42_im = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  regsB_43_re = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  regsB_43_im = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  regsB_44_re = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  regsB_44_im = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  regsB_45_re = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  regsB_45_im = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  regsB_46_re = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  regsB_46_im = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  regsB_47_re = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  regsB_47_im = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  regsB_48_re = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  regsB_48_im = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  regsB_49_re = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  regsB_49_im = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  regsB_50_re = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  regsB_50_im = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  regsB_51_re = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  regsB_51_im = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  regsB_52_re = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  regsB_52_im = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  regsB_53_re = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  regsB_53_im = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  regsB_54_re = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  regsB_54_im = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  regsB_55_re = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  regsB_55_im = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  regsB_56_re = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  regsB_56_im = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  regsB_57_re = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  regsB_57_im = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  regsB_58_re = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  regsB_58_im = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  regsB_59_re = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  regsB_59_im = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  regsB_60_re = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  regsB_60_im = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  regsB_61_re = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  regsB_61_im = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  regsB_62_re = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  regsB_62_im = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  regsB_63_re = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  regsB_63_im = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  regsB_64_re = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  regsB_64_im = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  regsB_65_re = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  regsB_65_im = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  regsB_66_re = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  regsB_66_im = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  regsB_67_re = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  regsB_67_im = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  regsB_68_re = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  regsB_68_im = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  regsB_69_re = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  regsB_69_im = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  regsB_70_re = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  regsB_70_im = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  regsB_71_re = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  regsB_71_im = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  regsB_72_re = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  regsB_72_im = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  regsB_73_re = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  regsB_73_im = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  regsB_74_re = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  regsB_74_im = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  regsB_75_re = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  regsB_75_im = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  regsB_76_re = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  regsB_76_im = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  regsB_77_re = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  regsB_77_im = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  regsB_78_re = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  regsB_78_im = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  regsB_79_re = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  regsB_79_im = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  regsB_80_re = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  regsB_80_im = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  regsB_81_re = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  regsB_81_im = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  regsB_82_re = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  regsB_82_im = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  regsB_83_re = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  regsB_83_im = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  regsB_84_re = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  regsB_84_im = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  regsB_85_re = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  regsB_85_im = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  regsB_86_re = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  regsB_86_im = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  regsB_87_re = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  regsB_87_im = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  regsB_88_re = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  regsB_88_im = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  regsB_89_re = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  regsB_89_im = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  regsB_90_re = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  regsB_90_im = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  regsB_91_re = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  regsB_91_im = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  regsB_92_re = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  regsB_92_im = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  regsB_93_re = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  regsB_93_im = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  regsB_94_re = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  regsB_94_im = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  regsB_95_re = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  regsB_95_im = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  regsB_96_re = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  regsB_96_im = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  regsB_97_re = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  regsB_97_im = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  regsB_98_re = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  regsB_98_im = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  regsB_99_re = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  regsB_99_im = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  input_point = _RAND_400[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
