module matrix_transpose(
  input         clock,
  input         reset,
  input  [63:0] io_matrixIn_0_re,
  input  [63:0] io_matrixIn_0_im,
  input  [63:0] io_matrixIn_1_re,
  input  [63:0] io_matrixIn_1_im,
  input  [63:0] io_matrixIn_2_re,
  input  [63:0] io_matrixIn_2_im,
  input  [63:0] io_matrixIn_3_re,
  input  [63:0] io_matrixIn_3_im,
  input  [63:0] io_matrixIn_4_re,
  input  [63:0] io_matrixIn_4_im,
  input  [63:0] io_matrixIn_5_re,
  input  [63:0] io_matrixIn_5_im,
  input  [63:0] io_matrixIn_6_re,
  input  [63:0] io_matrixIn_6_im,
  input  [63:0] io_matrixIn_7_re,
  input  [63:0] io_matrixIn_7_im,
  input  [63:0] io_matrixIn_8_re,
  input  [63:0] io_matrixIn_8_im,
  input  [63:0] io_matrixIn_9_re,
  input  [63:0] io_matrixIn_9_im,
  input  [63:0] io_matrixIn_10_re,
  input  [63:0] io_matrixIn_10_im,
  input  [63:0] io_matrixIn_11_re,
  input  [63:0] io_matrixIn_11_im,
  input  [63:0] io_matrixIn_12_re,
  input  [63:0] io_matrixIn_12_im,
  input  [63:0] io_matrixIn_13_re,
  input  [63:0] io_matrixIn_13_im,
  input  [63:0] io_matrixIn_14_re,
  input  [63:0] io_matrixIn_14_im,
  input  [63:0] io_matrixIn_15_re,
  input  [63:0] io_matrixIn_15_im,
  input  [63:0] io_matrixIn_16_re,
  input  [63:0] io_matrixIn_16_im,
  input  [63:0] io_matrixIn_17_re,
  input  [63:0] io_matrixIn_17_im,
  input  [63:0] io_matrixIn_18_re,
  input  [63:0] io_matrixIn_18_im,
  input  [63:0] io_matrixIn_19_re,
  input  [63:0] io_matrixIn_19_im,
  input  [63:0] io_matrixIn_20_re,
  input  [63:0] io_matrixIn_20_im,
  input  [63:0] io_matrixIn_21_re,
  input  [63:0] io_matrixIn_21_im,
  input  [63:0] io_matrixIn_22_re,
  input  [63:0] io_matrixIn_22_im,
  input  [63:0] io_matrixIn_23_re,
  input  [63:0] io_matrixIn_23_im,
  input  [63:0] io_matrixIn_24_re,
  input  [63:0] io_matrixIn_24_im,
  input  [63:0] io_matrixIn_25_re,
  input  [63:0] io_matrixIn_25_im,
  input  [63:0] io_matrixIn_26_re,
  input  [63:0] io_matrixIn_26_im,
  input  [63:0] io_matrixIn_27_re,
  input  [63:0] io_matrixIn_27_im,
  input  [63:0] io_matrixIn_28_re,
  input  [63:0] io_matrixIn_28_im,
  input  [63:0] io_matrixIn_29_re,
  input  [63:0] io_matrixIn_29_im,
  input  [63:0] io_matrixIn_30_re,
  input  [63:0] io_matrixIn_30_im,
  input  [63:0] io_matrixIn_31_re,
  input  [63:0] io_matrixIn_31_im,
  input  [63:0] io_matrixIn_32_re,
  input  [63:0] io_matrixIn_32_im,
  input  [63:0] io_matrixIn_33_re,
  input  [63:0] io_matrixIn_33_im,
  input  [63:0] io_matrixIn_34_re,
  input  [63:0] io_matrixIn_34_im,
  input  [63:0] io_matrixIn_35_re,
  input  [63:0] io_matrixIn_35_im,
  input  [63:0] io_matrixIn_36_re,
  input  [63:0] io_matrixIn_36_im,
  input  [63:0] io_matrixIn_37_re,
  input  [63:0] io_matrixIn_37_im,
  input  [63:0] io_matrixIn_38_re,
  input  [63:0] io_matrixIn_38_im,
  input  [63:0] io_matrixIn_39_re,
  input  [63:0] io_matrixIn_39_im,
  input  [63:0] io_matrixIn_40_re,
  input  [63:0] io_matrixIn_40_im,
  input  [63:0] io_matrixIn_41_re,
  input  [63:0] io_matrixIn_41_im,
  input  [63:0] io_matrixIn_42_re,
  input  [63:0] io_matrixIn_42_im,
  input  [63:0] io_matrixIn_43_re,
  input  [63:0] io_matrixIn_43_im,
  input  [63:0] io_matrixIn_44_re,
  input  [63:0] io_matrixIn_44_im,
  input  [63:0] io_matrixIn_45_re,
  input  [63:0] io_matrixIn_45_im,
  input  [63:0] io_matrixIn_46_re,
  input  [63:0] io_matrixIn_46_im,
  input  [63:0] io_matrixIn_47_re,
  input  [63:0] io_matrixIn_47_im,
  input  [63:0] io_matrixIn_48_re,
  input  [63:0] io_matrixIn_48_im,
  input  [63:0] io_matrixIn_49_re,
  input  [63:0] io_matrixIn_49_im,
  input  [63:0] io_matrixIn_50_re,
  input  [63:0] io_matrixIn_50_im,
  input  [63:0] io_matrixIn_51_re,
  input  [63:0] io_matrixIn_51_im,
  input  [63:0] io_matrixIn_52_re,
  input  [63:0] io_matrixIn_52_im,
  input  [63:0] io_matrixIn_53_re,
  input  [63:0] io_matrixIn_53_im,
  input  [63:0] io_matrixIn_54_re,
  input  [63:0] io_matrixIn_54_im,
  input  [63:0] io_matrixIn_55_re,
  input  [63:0] io_matrixIn_55_im,
  input  [63:0] io_matrixIn_56_re,
  input  [63:0] io_matrixIn_56_im,
  input  [63:0] io_matrixIn_57_re,
  input  [63:0] io_matrixIn_57_im,
  input  [63:0] io_matrixIn_58_re,
  input  [63:0] io_matrixIn_58_im,
  input  [63:0] io_matrixIn_59_re,
  input  [63:0] io_matrixIn_59_im,
  input  [63:0] io_matrixIn_60_re,
  input  [63:0] io_matrixIn_60_im,
  input  [63:0] io_matrixIn_61_re,
  input  [63:0] io_matrixIn_61_im,
  input  [63:0] io_matrixIn_62_re,
  input  [63:0] io_matrixIn_62_im,
  input  [63:0] io_matrixIn_63_re,
  input  [63:0] io_matrixIn_63_im,
  input  [63:0] io_matrixIn_64_re,
  input  [63:0] io_matrixIn_64_im,
  input  [63:0] io_matrixIn_65_re,
  input  [63:0] io_matrixIn_65_im,
  input  [63:0] io_matrixIn_66_re,
  input  [63:0] io_matrixIn_66_im,
  input  [63:0] io_matrixIn_67_re,
  input  [63:0] io_matrixIn_67_im,
  input  [63:0] io_matrixIn_68_re,
  input  [63:0] io_matrixIn_68_im,
  input  [63:0] io_matrixIn_69_re,
  input  [63:0] io_matrixIn_69_im,
  input  [63:0] io_matrixIn_70_re,
  input  [63:0] io_matrixIn_70_im,
  input  [63:0] io_matrixIn_71_re,
  input  [63:0] io_matrixIn_71_im,
  input  [63:0] io_matrixIn_72_re,
  input  [63:0] io_matrixIn_72_im,
  input  [63:0] io_matrixIn_73_re,
  input  [63:0] io_matrixIn_73_im,
  input  [63:0] io_matrixIn_74_re,
  input  [63:0] io_matrixIn_74_im,
  input  [63:0] io_matrixIn_75_re,
  input  [63:0] io_matrixIn_75_im,
  input  [63:0] io_matrixIn_76_re,
  input  [63:0] io_matrixIn_76_im,
  input  [63:0] io_matrixIn_77_re,
  input  [63:0] io_matrixIn_77_im,
  input  [63:0] io_matrixIn_78_re,
  input  [63:0] io_matrixIn_78_im,
  input  [63:0] io_matrixIn_79_re,
  input  [63:0] io_matrixIn_79_im,
  input  [63:0] io_matrixIn_80_re,
  input  [63:0] io_matrixIn_80_im,
  input  [63:0] io_matrixIn_81_re,
  input  [63:0] io_matrixIn_81_im,
  input  [63:0] io_matrixIn_82_re,
  input  [63:0] io_matrixIn_82_im,
  input  [63:0] io_matrixIn_83_re,
  input  [63:0] io_matrixIn_83_im,
  input  [63:0] io_matrixIn_84_re,
  input  [63:0] io_matrixIn_84_im,
  input  [63:0] io_matrixIn_85_re,
  input  [63:0] io_matrixIn_85_im,
  input  [63:0] io_matrixIn_86_re,
  input  [63:0] io_matrixIn_86_im,
  input  [63:0] io_matrixIn_87_re,
  input  [63:0] io_matrixIn_87_im,
  input  [63:0] io_matrixIn_88_re,
  input  [63:0] io_matrixIn_88_im,
  input  [63:0] io_matrixIn_89_re,
  input  [63:0] io_matrixIn_89_im,
  input  [63:0] io_matrixIn_90_re,
  input  [63:0] io_matrixIn_90_im,
  input  [63:0] io_matrixIn_91_re,
  input  [63:0] io_matrixIn_91_im,
  input  [63:0] io_matrixIn_92_re,
  input  [63:0] io_matrixIn_92_im,
  input  [63:0] io_matrixIn_93_re,
  input  [63:0] io_matrixIn_93_im,
  input  [63:0] io_matrixIn_94_re,
  input  [63:0] io_matrixIn_94_im,
  input  [63:0] io_matrixIn_95_re,
  input  [63:0] io_matrixIn_95_im,
  input  [63:0] io_matrixIn_96_re,
  input  [63:0] io_matrixIn_96_im,
  input  [63:0] io_matrixIn_97_re,
  input  [63:0] io_matrixIn_97_im,
  input  [63:0] io_matrixIn_98_re,
  input  [63:0] io_matrixIn_98_im,
  input  [63:0] io_matrixIn_99_re,
  input  [63:0] io_matrixIn_99_im,
  output [63:0] io_matrixOut_0_re,
  output [63:0] io_matrixOut_0_im,
  output [63:0] io_matrixOut_1_re,
  output [63:0] io_matrixOut_1_im,
  output [63:0] io_matrixOut_2_re,
  output [63:0] io_matrixOut_2_im,
  output [63:0] io_matrixOut_3_re,
  output [63:0] io_matrixOut_3_im,
  output [63:0] io_matrixOut_4_re,
  output [63:0] io_matrixOut_4_im,
  output [63:0] io_matrixOut_5_re,
  output [63:0] io_matrixOut_5_im,
  output [63:0] io_matrixOut_6_re,
  output [63:0] io_matrixOut_6_im,
  output [63:0] io_matrixOut_7_re,
  output [63:0] io_matrixOut_7_im,
  output [63:0] io_matrixOut_8_re,
  output [63:0] io_matrixOut_8_im,
  output [63:0] io_matrixOut_9_re,
  output [63:0] io_matrixOut_9_im,
  output [63:0] io_matrixOut_10_re,
  output [63:0] io_matrixOut_10_im,
  output [63:0] io_matrixOut_11_re,
  output [63:0] io_matrixOut_11_im,
  output [63:0] io_matrixOut_12_re,
  output [63:0] io_matrixOut_12_im,
  output [63:0] io_matrixOut_13_re,
  output [63:0] io_matrixOut_13_im,
  output [63:0] io_matrixOut_14_re,
  output [63:0] io_matrixOut_14_im,
  output [63:0] io_matrixOut_15_re,
  output [63:0] io_matrixOut_15_im,
  output [63:0] io_matrixOut_16_re,
  output [63:0] io_matrixOut_16_im,
  output [63:0] io_matrixOut_17_re,
  output [63:0] io_matrixOut_17_im,
  output [63:0] io_matrixOut_18_re,
  output [63:0] io_matrixOut_18_im,
  output [63:0] io_matrixOut_19_re,
  output [63:0] io_matrixOut_19_im,
  output [63:0] io_matrixOut_20_re,
  output [63:0] io_matrixOut_20_im,
  output [63:0] io_matrixOut_21_re,
  output [63:0] io_matrixOut_21_im,
  output [63:0] io_matrixOut_22_re,
  output [63:0] io_matrixOut_22_im,
  output [63:0] io_matrixOut_23_re,
  output [63:0] io_matrixOut_23_im,
  output [63:0] io_matrixOut_24_re,
  output [63:0] io_matrixOut_24_im,
  output [63:0] io_matrixOut_25_re,
  output [63:0] io_matrixOut_25_im,
  output [63:0] io_matrixOut_26_re,
  output [63:0] io_matrixOut_26_im,
  output [63:0] io_matrixOut_27_re,
  output [63:0] io_matrixOut_27_im,
  output [63:0] io_matrixOut_28_re,
  output [63:0] io_matrixOut_28_im,
  output [63:0] io_matrixOut_29_re,
  output [63:0] io_matrixOut_29_im,
  output [63:0] io_matrixOut_30_re,
  output [63:0] io_matrixOut_30_im,
  output [63:0] io_matrixOut_31_re,
  output [63:0] io_matrixOut_31_im,
  output [63:0] io_matrixOut_32_re,
  output [63:0] io_matrixOut_32_im,
  output [63:0] io_matrixOut_33_re,
  output [63:0] io_matrixOut_33_im,
  output [63:0] io_matrixOut_34_re,
  output [63:0] io_matrixOut_34_im,
  output [63:0] io_matrixOut_35_re,
  output [63:0] io_matrixOut_35_im,
  output [63:0] io_matrixOut_36_re,
  output [63:0] io_matrixOut_36_im,
  output [63:0] io_matrixOut_37_re,
  output [63:0] io_matrixOut_37_im,
  output [63:0] io_matrixOut_38_re,
  output [63:0] io_matrixOut_38_im,
  output [63:0] io_matrixOut_39_re,
  output [63:0] io_matrixOut_39_im,
  output [63:0] io_matrixOut_40_re,
  output [63:0] io_matrixOut_40_im,
  output [63:0] io_matrixOut_41_re,
  output [63:0] io_matrixOut_41_im,
  output [63:0] io_matrixOut_42_re,
  output [63:0] io_matrixOut_42_im,
  output [63:0] io_matrixOut_43_re,
  output [63:0] io_matrixOut_43_im,
  output [63:0] io_matrixOut_44_re,
  output [63:0] io_matrixOut_44_im,
  output [63:0] io_matrixOut_45_re,
  output [63:0] io_matrixOut_45_im,
  output [63:0] io_matrixOut_46_re,
  output [63:0] io_matrixOut_46_im,
  output [63:0] io_matrixOut_47_re,
  output [63:0] io_matrixOut_47_im,
  output [63:0] io_matrixOut_48_re,
  output [63:0] io_matrixOut_48_im,
  output [63:0] io_matrixOut_49_re,
  output [63:0] io_matrixOut_49_im,
  output [63:0] io_matrixOut_50_re,
  output [63:0] io_matrixOut_50_im,
  output [63:0] io_matrixOut_51_re,
  output [63:0] io_matrixOut_51_im,
  output [63:0] io_matrixOut_52_re,
  output [63:0] io_matrixOut_52_im,
  output [63:0] io_matrixOut_53_re,
  output [63:0] io_matrixOut_53_im,
  output [63:0] io_matrixOut_54_re,
  output [63:0] io_matrixOut_54_im,
  output [63:0] io_matrixOut_55_re,
  output [63:0] io_matrixOut_55_im,
  output [63:0] io_matrixOut_56_re,
  output [63:0] io_matrixOut_56_im,
  output [63:0] io_matrixOut_57_re,
  output [63:0] io_matrixOut_57_im,
  output [63:0] io_matrixOut_58_re,
  output [63:0] io_matrixOut_58_im,
  output [63:0] io_matrixOut_59_re,
  output [63:0] io_matrixOut_59_im,
  output [63:0] io_matrixOut_60_re,
  output [63:0] io_matrixOut_60_im,
  output [63:0] io_matrixOut_61_re,
  output [63:0] io_matrixOut_61_im,
  output [63:0] io_matrixOut_62_re,
  output [63:0] io_matrixOut_62_im,
  output [63:0] io_matrixOut_63_re,
  output [63:0] io_matrixOut_63_im,
  output [63:0] io_matrixOut_64_re,
  output [63:0] io_matrixOut_64_im,
  output [63:0] io_matrixOut_65_re,
  output [63:0] io_matrixOut_65_im,
  output [63:0] io_matrixOut_66_re,
  output [63:0] io_matrixOut_66_im,
  output [63:0] io_matrixOut_67_re,
  output [63:0] io_matrixOut_67_im,
  output [63:0] io_matrixOut_68_re,
  output [63:0] io_matrixOut_68_im,
  output [63:0] io_matrixOut_69_re,
  output [63:0] io_matrixOut_69_im,
  output [63:0] io_matrixOut_70_re,
  output [63:0] io_matrixOut_70_im,
  output [63:0] io_matrixOut_71_re,
  output [63:0] io_matrixOut_71_im,
  output [63:0] io_matrixOut_72_re,
  output [63:0] io_matrixOut_72_im,
  output [63:0] io_matrixOut_73_re,
  output [63:0] io_matrixOut_73_im,
  output [63:0] io_matrixOut_74_re,
  output [63:0] io_matrixOut_74_im,
  output [63:0] io_matrixOut_75_re,
  output [63:0] io_matrixOut_75_im,
  output [63:0] io_matrixOut_76_re,
  output [63:0] io_matrixOut_76_im,
  output [63:0] io_matrixOut_77_re,
  output [63:0] io_matrixOut_77_im,
  output [63:0] io_matrixOut_78_re,
  output [63:0] io_matrixOut_78_im,
  output [63:0] io_matrixOut_79_re,
  output [63:0] io_matrixOut_79_im,
  output [63:0] io_matrixOut_80_re,
  output [63:0] io_matrixOut_80_im,
  output [63:0] io_matrixOut_81_re,
  output [63:0] io_matrixOut_81_im,
  output [63:0] io_matrixOut_82_re,
  output [63:0] io_matrixOut_82_im,
  output [63:0] io_matrixOut_83_re,
  output [63:0] io_matrixOut_83_im,
  output [63:0] io_matrixOut_84_re,
  output [63:0] io_matrixOut_84_im,
  output [63:0] io_matrixOut_85_re,
  output [63:0] io_matrixOut_85_im,
  output [63:0] io_matrixOut_86_re,
  output [63:0] io_matrixOut_86_im,
  output [63:0] io_matrixOut_87_re,
  output [63:0] io_matrixOut_87_im,
  output [63:0] io_matrixOut_88_re,
  output [63:0] io_matrixOut_88_im,
  output [63:0] io_matrixOut_89_re,
  output [63:0] io_matrixOut_89_im,
  output [63:0] io_matrixOut_90_re,
  output [63:0] io_matrixOut_90_im,
  output [63:0] io_matrixOut_91_re,
  output [63:0] io_matrixOut_91_im,
  output [63:0] io_matrixOut_92_re,
  output [63:0] io_matrixOut_92_im,
  output [63:0] io_matrixOut_93_re,
  output [63:0] io_matrixOut_93_im,
  output [63:0] io_matrixOut_94_re,
  output [63:0] io_matrixOut_94_im,
  output [63:0] io_matrixOut_95_re,
  output [63:0] io_matrixOut_95_im,
  output [63:0] io_matrixOut_96_re,
  output [63:0] io_matrixOut_96_im,
  output [63:0] io_matrixOut_97_re,
  output [63:0] io_matrixOut_97_im,
  output [63:0] io_matrixOut_98_re,
  output [63:0] io_matrixOut_98_im,
  output [63:0] io_matrixOut_99_re,
  output [63:0] io_matrixOut_99_im
);
  assign io_matrixOut_0_re = io_matrixIn_0_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_0_im = io_matrixIn_0_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_1_re = io_matrixIn_10_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_1_im = io_matrixIn_10_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_2_re = io_matrixIn_20_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_2_im = io_matrixIn_20_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_3_re = io_matrixIn_30_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_3_im = io_matrixIn_30_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_4_re = io_matrixIn_40_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_4_im = io_matrixIn_40_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_5_re = io_matrixIn_50_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_5_im = io_matrixIn_50_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_6_re = io_matrixIn_60_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_6_im = io_matrixIn_60_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_7_re = io_matrixIn_70_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_7_im = io_matrixIn_70_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_8_re = io_matrixIn_80_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_8_im = io_matrixIn_80_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_9_re = io_matrixIn_90_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_9_im = io_matrixIn_90_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_10_re = io_matrixIn_1_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_10_im = io_matrixIn_1_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_11_re = io_matrixIn_11_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_11_im = io_matrixIn_11_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_12_re = io_matrixIn_21_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_12_im = io_matrixIn_21_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_13_re = io_matrixIn_31_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_13_im = io_matrixIn_31_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_14_re = io_matrixIn_41_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_14_im = io_matrixIn_41_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_15_re = io_matrixIn_51_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_15_im = io_matrixIn_51_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_16_re = io_matrixIn_61_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_16_im = io_matrixIn_61_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_17_re = io_matrixIn_71_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_17_im = io_matrixIn_71_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_18_re = io_matrixIn_81_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_18_im = io_matrixIn_81_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_19_re = io_matrixIn_91_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_19_im = io_matrixIn_91_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_20_re = io_matrixIn_2_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_20_im = io_matrixIn_2_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_21_re = io_matrixIn_12_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_21_im = io_matrixIn_12_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_22_re = io_matrixIn_22_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_22_im = io_matrixIn_22_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_23_re = io_matrixIn_32_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_23_im = io_matrixIn_32_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_24_re = io_matrixIn_42_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_24_im = io_matrixIn_42_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_25_re = io_matrixIn_52_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_25_im = io_matrixIn_52_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_26_re = io_matrixIn_62_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_26_im = io_matrixIn_62_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_27_re = io_matrixIn_72_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_27_im = io_matrixIn_72_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_28_re = io_matrixIn_82_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_28_im = io_matrixIn_82_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_29_re = io_matrixIn_92_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_29_im = io_matrixIn_92_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_30_re = io_matrixIn_3_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_30_im = io_matrixIn_3_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_31_re = io_matrixIn_13_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_31_im = io_matrixIn_13_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_32_re = io_matrixIn_23_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_32_im = io_matrixIn_23_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_33_re = io_matrixIn_33_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_33_im = io_matrixIn_33_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_34_re = io_matrixIn_43_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_34_im = io_matrixIn_43_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_35_re = io_matrixIn_53_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_35_im = io_matrixIn_53_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_36_re = io_matrixIn_63_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_36_im = io_matrixIn_63_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_37_re = io_matrixIn_73_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_37_im = io_matrixIn_73_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_38_re = io_matrixIn_83_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_38_im = io_matrixIn_83_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_39_re = io_matrixIn_93_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_39_im = io_matrixIn_93_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_40_re = io_matrixIn_4_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_40_im = io_matrixIn_4_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_41_re = io_matrixIn_14_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_41_im = io_matrixIn_14_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_42_re = io_matrixIn_24_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_42_im = io_matrixIn_24_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_43_re = io_matrixIn_34_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_43_im = io_matrixIn_34_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_44_re = io_matrixIn_44_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_44_im = io_matrixIn_44_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_45_re = io_matrixIn_54_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_45_im = io_matrixIn_54_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_46_re = io_matrixIn_64_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_46_im = io_matrixIn_64_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_47_re = io_matrixIn_74_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_47_im = io_matrixIn_74_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_48_re = io_matrixIn_84_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_48_im = io_matrixIn_84_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_49_re = io_matrixIn_94_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_49_im = io_matrixIn_94_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_50_re = io_matrixIn_5_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_50_im = io_matrixIn_5_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_51_re = io_matrixIn_15_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_51_im = io_matrixIn_15_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_52_re = io_matrixIn_25_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_52_im = io_matrixIn_25_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_53_re = io_matrixIn_35_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_53_im = io_matrixIn_35_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_54_re = io_matrixIn_45_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_54_im = io_matrixIn_45_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_55_re = io_matrixIn_55_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_55_im = io_matrixIn_55_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_56_re = io_matrixIn_65_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_56_im = io_matrixIn_65_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_57_re = io_matrixIn_75_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_57_im = io_matrixIn_75_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_58_re = io_matrixIn_85_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_58_im = io_matrixIn_85_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_59_re = io_matrixIn_95_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_59_im = io_matrixIn_95_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_60_re = io_matrixIn_6_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_60_im = io_matrixIn_6_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_61_re = io_matrixIn_16_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_61_im = io_matrixIn_16_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_62_re = io_matrixIn_26_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_62_im = io_matrixIn_26_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_63_re = io_matrixIn_36_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_63_im = io_matrixIn_36_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_64_re = io_matrixIn_46_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_64_im = io_matrixIn_46_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_65_re = io_matrixIn_56_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_65_im = io_matrixIn_56_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_66_re = io_matrixIn_66_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_66_im = io_matrixIn_66_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_67_re = io_matrixIn_76_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_67_im = io_matrixIn_76_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_68_re = io_matrixIn_86_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_68_im = io_matrixIn_86_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_69_re = io_matrixIn_96_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_69_im = io_matrixIn_96_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_70_re = io_matrixIn_7_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_70_im = io_matrixIn_7_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_71_re = io_matrixIn_17_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_71_im = io_matrixIn_17_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_72_re = io_matrixIn_27_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_72_im = io_matrixIn_27_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_73_re = io_matrixIn_37_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_73_im = io_matrixIn_37_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_74_re = io_matrixIn_47_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_74_im = io_matrixIn_47_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_75_re = io_matrixIn_57_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_75_im = io_matrixIn_57_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_76_re = io_matrixIn_67_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_76_im = io_matrixIn_67_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_77_re = io_matrixIn_77_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_77_im = io_matrixIn_77_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_78_re = io_matrixIn_87_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_78_im = io_matrixIn_87_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_79_re = io_matrixIn_97_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_79_im = io_matrixIn_97_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_80_re = io_matrixIn_8_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_80_im = io_matrixIn_8_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_81_re = io_matrixIn_18_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_81_im = io_matrixIn_18_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_82_re = io_matrixIn_28_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_82_im = io_matrixIn_28_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_83_re = io_matrixIn_38_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_83_im = io_matrixIn_38_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_84_re = io_matrixIn_48_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_84_im = io_matrixIn_48_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_85_re = io_matrixIn_58_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_85_im = io_matrixIn_58_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_86_re = io_matrixIn_68_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_86_im = io_matrixIn_68_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_87_re = io_matrixIn_78_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_87_im = io_matrixIn_78_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_88_re = io_matrixIn_88_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_88_im = io_matrixIn_88_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_89_re = io_matrixIn_98_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_89_im = io_matrixIn_98_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_90_re = io_matrixIn_9_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_90_im = io_matrixIn_9_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_91_re = io_matrixIn_19_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_91_im = io_matrixIn_19_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_92_re = io_matrixIn_29_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_92_im = io_matrixIn_29_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_93_re = io_matrixIn_39_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_93_im = io_matrixIn_39_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_94_re = io_matrixIn_49_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_94_im = io_matrixIn_49_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_95_re = io_matrixIn_59_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_95_im = io_matrixIn_59_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_96_re = io_matrixIn_69_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_96_im = io_matrixIn_69_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_97_re = io_matrixIn_79_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_97_im = io_matrixIn_79_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_98_re = io_matrixIn_89_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_98_im = io_matrixIn_89_im; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_99_re = io_matrixIn_99_re; // @[Matrix_Transpose.scala 22:31]
  assign io_matrixOut_99_im = io_matrixIn_99_im; // @[Matrix_Transpose.scala 22:31]
endmodule
